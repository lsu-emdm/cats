BZh91AY&SY�|�y�8߀rx����� ����ay�       } M�Fd����H: C�6�G
��Q�U]�Ю	��h�.�`:       
            �� "(R� (U( ����T��U)Jf         =�   � -�=�x
=���X�ٸ�;=��8n)�o/N{u�F^�:pJ�rb�]�ǀ	y�R�
`�(�8 ��n���`)�wu��x�T�w3�����)N�t(��p� $\   q� ���e��-�gϾ�o�x�}�������j�3�Ӽ�/Z��u}���\�����j���}G��s�{j������@0�Z���x�v���
��ꗽ��ں��=z�y�z��|�}j��Gp��o}j�����۷���k�UW(�    �   8<}U�}�>�_}}��}����=�M����q�}�6�ή��q�m�=���x��]�=�m.Z�m�7^� wo.G�/z���U�o�����}�܅��^}o��|�������}o��k����>��z��W�<|   �
� <���z/�v�^�{�����}{�[��&�ן |��|e�|f��wof�w{7�����x���M�7}����9|�O=��|�K�]�Խ�z�����|Ǖn��8s���������{ֲ������`w� �|   �O@ �<)�}�suJ�n�m^�;���|܋��U�^Ǽ��5<��͹g�����m�<t���%����O6�� 6_w�ﯽ�p<R]��y�ﯮ^l�=���:�[���f��.�ٞ���/{w�kũ|۾n��� @        
�jR�Q�       i��)J���&�@ ����z�R<�D@`���2MMjy�"����ɠ @  S��I��J�M !�4i�F  B��J@Ц��C&�='��CF�MM1)��?t��������ǯ��X{{}�^��UEW�Ռp��������� ����@U]?�**��7�_������/��������?�߿�����)=TUb�tl�* �nl�z`���?~`u����'��罚T�(�����o��.�џ���������V�h@�C�%Pu*��R���L���r�V�ZQDh�C�u(�@P�� jD(P�QJ � ���
���T5 (P��U�T浤V����Di�$]k\�"��]B�
*4�
ЮJ�@d�PH�"9*�"�	�
' @Ԣ��Au"��AhG$��R�B�V�R :�B��J��]@�U�+�� )B�%C����%PiS!\�JE�b*rh �]ku�Ew"�*��T5(�jU�(С�Ap�Aܛ�&��3 ��r:��Z5n �r��4!�+�n
�7	�5�5d��5<�7+Bj!i���
nC#�P�BP�NG$��17��:�&��%��r7�Rd!JR���<���(P
��L�	2ZrJ�#q��.IBd�&�IAIo䦳# 0� r
9.��ԉZ�.�)���rL�
i2A���7nH#�h
MC�y!�b��Լ���u	�Mș���a�P9)Bji��C%(�ZS������w�kr.�CR�B���%�2�rP��)!�i)
������i2E2)ԙ �D��7@:����䁻q�Cr����5���7��@��	31FC�5N�&� u��Y�9Re�d�6`�Rd�%!AK��rGR��V��
���%\�5 �kVb9K��-��`��K�!�nu+���a���ug0r9d!���)y.��@P)AA�7!��p�ʗ$)rirV����((hZA�������2
 )���r5% ��A��Hjە��H��Ժ�hu	�u dJrP�T�Gp9�R�.Y P@�P���!J�@�H�H�B�(�
Ү��P� ;��G%DhP�V�ZT�F� ���<�g�����x������.���b&�)��u&Ǧ���[YK�x0�[����}�V��ʩ>v�ܻ-��c��̔AN�
���s+�yoQ���=U�͝|������b�v�v��)�=^E�_�=T(�y�up�.תZK���[��Fk�yTĩy�]�:.�lb�1���z���-�^e�*���%�T�
�o:�s^�xUpF(UMD@�f(g�+������������[b�ר�؟<�Su�=���3ua�S1{���<�ne>��L�lNX���U��j��W�}ֿe�ޥm�K�\�\�%���I���H[j	��$I�N���e�v��
��r:�Zys\y���[�gG'�p8\����#3��'	����'I8͌�&�q�'ܫ޶�!P��xSZ��</0��T)�{�6�v��U�V�z��"P�R��,kZ�fu)Uk��Y���:�S%+^ŊЭjh�SV���n:ۅI�!:���Z�-�c3��Tֽ�p�E)I	�L�����y业�Ovo����vpcZy���A���6p�"�]���΋�<��'�������!)q�}|;6��;�Y���o����B��l�L0�>{����^�[�^J%;�BPK)JN��R�k�rj�/���s��H�x_=}����avy,}��y͈�󽯓{	�o&�
�;����F.�ai��������N�3���vk:#Fl�G4WK�q��mѻ���:�\ѯy���ב	'Y
e��d��J���ZM�X�犈ʟ<����ʬ��Je�2!2.s{�~��W � ��m��Q�͜9��/5�P����x��:�]�%�����3:a�<�"��gk�D�*i���iR�zt�5VsU�٣�A��w	Jw	�&Bj��2P�%Bj��%	Bd&Bu	Jjp�'P�&BP�%	��'p�&�2���:��P�BP���:��ٛ������,G~j������=����K�Mi�ddl�ѽ���q:#�c����h�yv����5NI���m�\w��<�'r�%	��	����!(L��2!=�́��%	BVs�Aqu�QZ���&�&�_%�'��9���5Џ`:x�3��nv��y�8��o#X]�v�X�f��;+'���{w���F{�Y�4xm�΋]֍�$�F������d�y�1�1e��7=���&�o���w�E؜�h���:�M�N��<���Ѣ;4�n\|��a;�T�wa����>^�|�ga��>Ád�js����vO�܄{o'i=��9�q���7�����Ra��7	Bd�	�M�PWo{�_�0����e�g:#[��Xlۇ�p21Ŝ�v��5��l��̚İ�w:+���qd�o���y�ǐa�uJ�T++ɆN�B��k��H|���O[�\7	Br�J��)J�L��(J�J!)J�MBP��m�sC��+���t�b'����&�2��)M�P���L��2��)N�(J�N�2P���M�r�MBP�	BP�%	����(Oa2������J��%	��&�2��	�J��=��(J��(J��J!(MBd�	��	��%	����MJP�	�M�d&�2�J�=�|/;��B�ӳpc�{甴4�>w(x�xB�Hg�%�R��(=�b�V�L����w@
�%�4�W����Hg��EZ��y[�c@̨IBd%	I;.	Ny�Q�2-���rLj��!��iw�Kqu	Jr��J!2!5	�%=�Z�}$��#�@09Jg)�er��*nK��9�L��,g�f��@����P�eBj���Թ՚���5���g-oC��ц���>�;��(O!2S��%	��%	BP�p�ɹ�R�b�F��ҴPP�� �HJGH�uA8�B��Y=��i�����<<͒G�G`2X����ړ n�������ý��v�l��C��X�w�	��\���C��&������w�x�d'p������t��ܧ!(J���z�G~.�Ȟ@dD]`<�;��y�	C��Lߤ�F��(�!C(�%�/5��+վ�YW�V$��]��y�HA
EP���J���!=�;4;�;t�w�}���=�Ѓ�)^���r�v�eO O#8^b0�=���|䞺CO&���n��᛻;I�!�	5�K�}{�B�{n����J��LD+Y4����
��fL���JD
���7HO'ɡ�:�{���yf�i]ïb����&�FS�Զ()%	Bu	Jj�J�M�P�	�MBR����L��j�g�K�GD�PO����yo1�#̌,^3nKՕ>1��z��t��_=�F��^�3<(%=+Kq��@�l�G;:<N�Q�=vu�x���7�ߕ��<��(v�E����:O+�G|��Ѿ=w׹��掍y���12t���aky�V��r�ѷ}��p3{7`N���;�j�]jt�Ɯ��gl�ou�쎖e�#��Fj7�Z8�Fe<8n�SV�e�ݽp�o�3���f��vl�<�B�
&�!E{�k�J�����C2��ߩ������4�2��ͩi����Sc;(P3;<*M����F�d�!���+G���/kVe�SSs�E5#��%z��񞌱�Ox g]�����e��ST$��,��|�8�������&*B�BԞ%
j	eW^��45	��+�I�3����]��&q�	�������Q�=�����ö7�)�F�������3 ���A�͉\M��Ѵ�d�3ud/av����Y�-�c;B�s���^<\���%&�!(�ѳq���8F�bY	A�r�ѐd��%bA�	I��K�A����+
�6�xa���ָf��%c�N�������3���S��1RhNd��h�F��s��y{�xh������Ŭ�;����l�{�Od�)�i�;.}�=���k^�w���F��nyY�>�ٹf)#;�՗��gi=���f������xNn;��,ﱞ���%����zN�N�8���L�<�����gi��U{��~i���}x͸�RD�|MV�z)��y�[ho0��J�Lŉ��%*Ry�y)8Db���+2S��ОS�+X�yPԐ�B���g�c�U	:P��/V��7�U�j��Z�^g[��5�K|����Ӯ�k|��ٷ��$�2ӱՁ�e��ox��MÃ	��y�8Y7�Ӭ󝤗�(���{�7��������g��,�"D�ﳒ١ӵ�s�WI���k���os�:4[�G<��B�Uv_Z��bN��pI%�{��.9	BD8c�9�Hd�e�D�@d8hԞ�5��e���c�5��Lc#C	BS�dh�F�[04��p�+Hd;�O5	BR���5��ߤַ�@׌�Xhݚ���˫^i���۬�hN��{N1�ÞƓ�����E���7'F��=w��;{w<�E�A�y�z�Gg]�wh�#�.�i��ٳǣ\��zQsf�.���Z�9��N�@�}BŃ�̨����8����^���A�VT�?��G��N�I���j_)3�s�v��r�k�u�۹��Qϭ��8�{���#��D<��)�=>�YpE�y2%74bz��>��Θ{��7�N��SO]C_b�a�:�y�v� ��A�H��������"�v��")�K"�}eڎ�e�'�Y!Oy��~�S�hX�&#!:�u0�U�[]��웇R�U������S�nay�zɿW�U�P�QsB�=������-4܍��Yo�ճ]-3�-����Me�
��lif��"Pب�\�n���V���k�\��,/,��WFY�ml�$��D�Y�l�S���Zi1��2�Ka�K+]�o4�R�7��7��
��Y�-T��4�fa�䱶���ܶWr�]�ˬ�[�Y�n$��d�]�m�-�`��氶�Cl�G@�S;�{��~���������������g�����~~l�j���y�#���D��*�m�%��                                          ��                                                                    	                         Pz               h      -�H                               ~�                                                                          �   �  -�                  �=        �        �z                                                ��ph�3B�٥Z��af�[mq��[�lq�m         �           �              ��     v�               �  �          �m��  �` 2   n�  �           އ�           �            R�            �         �@ �  ��        )@    p    �    ��         `        C� �     )@      @     �   ���        �-�        �            R�    հ �p 9  �J  d ��  ��� )@A����� �p �@
P`8 p (0 8��  �J  d �� 2 R���� )@A����� �p �Cѐ�  �J  d � � (0 8��                                       C�                             p          H                        m  �z     	  �q�2m����䎵�%����5�&�`                  �   ��                                                    ��                  [@       ����������h~�����f��m�Wb�� Me�$ڶ �ɶ׫m�j�p��&�Wn��w7W.�-�m�V��Km�2����fH�p0t�颬4c-	�J�Ȋ�" $��.F �PZ�����[v1�(�en���&shڠ�8�0�#L���cWK:��MoZj���W-H6��N���N�g[m��&݅�Qe�e��-�b����X�ѕ����*�,A�U� 	UT� n�
P ��pڐ[m�� 8�@ ���j̺�඀� ��#v�cN�m���m�� /Zm������[�m��� m�f�,�c� $�|��c��۶�m� @����v p8v�ێm[�  ݶ$mY�Zl��I��e����[t�8�R��k [Kd�2 6�  'R�:]��׽�Y@���kH�T�P�l��ʬݳ�#��]e�Q ��ٍ�]kde�M���c���Cm� ���M9��%���V�%� V�$��k`N�jڐkFF�֛u�Cm�� ��uM�Z�U]�qԱB�!�9u��7[4�t���m��:B�m����Z$�q�Y�ܶZ�ڃ���a ]������  8�:kt���h�0V�].|��H�R��^�lK.�]$K��m����b+�6�lǈ@�ca��lI Ht��W^ԡzd�  -�$I�Ŏt�լe�l\ɦ@"��,��4�������"E�T�    �#�b� 6� H   �n�[zې�t�1z�H[dK�d�@	 m�  ����m�[��� �K���d�۶�Ji䲂� p $ YKu��m8 q"ɺlo�k@k5�-�gڶ�6	�   m��m��A�D��h�-�d��cm6��	e�{��ؚ���-���&�-���n͵������\�]�ѠF����aˠ�J�i�EP���mrΐ6�m�Iz�A#GP��β.����q$�2�&�F�y���פ���9���# �"��A�U��81]��i�z��׬^p䅶C���P�JBh U�6��n��;k�-�@�����-�v�i��-�u� �hk%��2wH�  ���H@R �d\������m�J�;n�6�ۣ\�  ��f+����wL�k�m'I�9�m{M� mI�w�-��� �6F���[�6�:�HmѬ�  �mmH�I�m�m��fM� z�-��nUtŴ�,6�hM@6�ml8���6#m-�6�[%���8�g   m����۶�E�պ� ;Z���Y�mz�[m� ����� 	���n�6.�ڳmi��]5�@I��ۢ�d�[HM���mn�gKR�K�,�2�/���9Z�mr��N�l��'��ޡ]cp�$��m����mI#�$�ݳ�I'�w����r��f�Y�9m�|�n�Y)o�
���a�b+��X����Q.�pռʶklvߑ�oxC���i��<����度�&�dogm��Mz�9�_ m:,]�L[��z�:� S�lr�H̕˶ �6�������}���9��-�j�(�-�[�e3��J[1��^�e�h�Il���[h��Ckm֮(,�͙�F;V�1<x�m���-�혶��%�sm�-Ը�k��&M�٥�6���d䓥�,�f��ke��h�����P����"�k�,6�m�F��-�Z۶�Ɩ�B1CjFڬöbâ�V�
�d�Im��6ݷ�M��ז���g$qoSm�8H��jض�����'ڵ뀶�����`�n��݄�-$�&�ap�o�\�m� 6�agYJݨ x,i;l�N9e��f�*dL����f-&�Qڮ-e�M��K76E���f�+�H�`��i6�\ �Z� ��p�c�  ��l$u�M�u[U�M�IIo
Yn�  �;m�l��Iƺ�l����Z1vֺ�:�k� �l�6	Vb3lY@U�v�d.�T���h�kR�j�j�m4j��+�ji�6ܠc�ŭ�-�e�^�N�]�.֠Z6ͪ�[F�6V�Ѭ-���)XP��Dj�J��P��m�F��f�sK��@��Q�` m4�vV�ƪ�%�am�ر%�yl�Z�g\eٵT��f�ui�k���h*� v��m��-��D.�θ[A�l�9$�l-�t�m� ����	�[@�I@��D�n�gd1�iU�S0��B �q�kh���m�u�R�X��ɵ��Xa�bѵ�xf���6�b�4u��Y�MD�!mͤkn��h�]Z/[��ٙl�m4���J�[I������7)r݋l�l���M$�Z�v�j鬂8�΄�N�׷ny�lߟ�� *
������  �����������DT?����_�4dl�U�k3N�8�Z�d���Z�yA��Ѳ4���3q"I4��a]-���Y-y/9yt��ˡ"�Yt���s3�嘓NHʹYY&�5��09�GY!	��X9����?��TAz�@�ß���E_�� �pv�C��FC�	����JB`�@ t�'Jb�0�.�1Sai_ RQ�@�8��H��6�*Z���/�	��Bb�H�UX�)(tt��&�d"H�&c�t!�}U${C� ���P�HG�v����}F��CB`���wDT�22& b�2L�Bj�8�P�D1<{�S�Skؐ�Y��{TM�����0;�h�*J�P�e&WJ*�zJb�����x�8mS��c��#��WH���LA�N�I<#p�E3�����N�NhC���FG:^ �h�� i ���1��t� ,t*&�0��:�
�b�`,Tt t=��B��� \z�}�9A��)؞/�m#)��|�\Dz@]�R0b�H� K�GU�0^0�
H�.�_A�Б�i��U�i��آ�� ��lT������@�
��@�8*�lG���Cl���M���%�u������ X�?������e�/O������5Lş�Y�7k��hu�J��(J��(J��(J��(JR��(J��(J��(J��(J��*����)J��(J��(J��(J%�
��(J��(J`��(!�	���Ր�0T	HB�d�����@*�d*��"�T�A�A�A�A�A�A�A�A��R�h"JDhA+0DhEB����%	BP�&f	BP�%	BP�����ШШШШШС��(J��&3$�&��(J��(JBP����(J��(J���(J��(J��(L���(J��(J���(J��(J��(L���(J��(J���(J��(J��(L���(J��(JP����(J��(J���(J�Mf��(JHr��(�3�$�(J��(L���(J��(J���(J��$���(J��J��Ƅ�(L�d����J��KBP�%	BP�%	��P�%	BP�%	BP��%	BP�%	BP�%	��P�%	BP�%	BP��%	BP�%	HNBP�bE	BP�&f	BP�%2d%	C�P�%	Bf`�%	BP�%	BP�&f	BP�%	L	BP�%	��P���%	�f`��2��*BP`�%	BP�d��%	BP�%	Bf`�%	BP�%	BP�&f	BP�%	BP�%	Bk0Jr�U_�Y��3���
j�BM#�?}<�q�}6ߘ�v�       �            [@6�  8 m�   l     m�              6��   l p�i06�	       e��n��@     �m�l   � @H�8  m� 8       dl  x     m�	  6�a�   C�-�8���b  d �� 2 R���q@A� �m    ��      �    �mK.��\Ƞ  ���    p     �     8�5�"i�r��̗mt�*"���"+�#�U	)��,��
������d��Fl4@f̢W.�c���v�B+��#F����jͮ�@E�4jѡ����~��y4���s�dMl��V��i�!�ܬ]��˃M2M����ĥ�e����Z�(�BoO>{��oM���EB�Λ l�[6�4-�q��.0��pj�u����,��e�f�ɑ�f�m�{��^��Zj�n*B�����t�\[�f�k�Z]-F�Fb;�>���� ���b&�nV�8�Y����xyUK6��h �%]��+LM�c�
��,����f�]̴ֺh�L��!�H rJ#�/�2��C'UC��U���(���`�0͞�ֲ��q	���Ұ�]0�ڹu��m���-ͭ�Q�6�-��v��en��
��ǙTյ�&G��g���o�۵�j�M���j�m�э-�nԵ,~s�>�{�x;���1x,�^$@��)���4��6X�c;]~Bj�}7b�]�{_X��]콛�Q �*�����J�>�����8$��1D�ڌ
/E�	>E +*>�!��h	}g���C����U�W W�����Ο�@l m -�6�  -hI{M� �� �M�2pm� 0�cn؝	)E�2�� ����`�`[m�A1��kp� �rg�{��v��N���@W6�f�Xk3���ي��̸�����͙\pŗ@���ei����/�5��4�qBh�X���3�l�/j ��oˢM�)���������9�����Ns��C`50nS1m��bR�Yn��%�`��.źR륛���/�|��@݉��Ƞ=��z�y�G�P	�J����2�;qCw!P����v���u�!K��x���q�݆�̍�C���X/fmR���:����C��k�ͥ�ݖ�o��F?fW=��3$T�R5)B9-}��+���^=�\�}촼�{$���F������i�M͛�D^M�9�$p�l6���.��ʢL�RLB�D��W�n��7bw��K�슅�,�F�!���G$��ٔFd�53c&�Q�T�3e-�dm5����u��*10�{�Kۻ-���ѹ�ʕ���,}�C��#�D�7�vZ_�-t�et��{-w���|� ��U*p#���E�n°�ͥ�ݕ�^O��$���mr����YU p�sE����&.�na6T�E.؀#wg'{i�i�i-�0/g���؁]�m,��j<�ݨ=���9)iP�0����j�vR��wm�6v"�Nl�d��)MU(J����}߳,!QTPU����]���<��m�=yg�0�~ݩ5{^5D:����*%�3c��u��{v�&^��m/LS���CQ�Ik����{��h_fe�s�����߼�������+��r�Sck���.e�l���LF4n�$�r��;�:58�6�bX�P�ҡ�n�a�)z��K����|��L�*(9U%��̊�ן�-Y����{gi_�}yi�iNH��۴���O�$�z%�߷�_wJ�B��u�!K��x��X�݆��͵��-���*A�+ 2��<Ϟ˵�+�L����T�}�fZ�3"_w����6f�s>ܭ���F ��y-���t Svu��NΪ�@q)5^U�.�D����$"�SUJ��>���}�2׏fV�qS_}��Y��U5 �	T��Q/}��fL���k�d��̥"�<�I�x�8�%ɗ��Znl5߲l32Z���oc���6�(xJT"ba����3%-�nҔ��9�\��P��E*U��2.�R\�M��ݭ\:{�"�9���I$�  ��[Am    C[n� �e� $g@  ��$g��0g6�2 R�m�` -����[ݽ[v�������A����KU���51~c���Ԗ�R�溋l��W�b�c.��XD(Z�,l�\�մ����μK��y6)-7fڰ-�*�:�i���CA0y~wv��W���\N�����#;��j�
��Z5��[:i�m���o/*��e�C:��jU7�{]8��Dq�I\�AQR�4��nב���߲U�d����B�wP�9h3v>d�0��ؕ�ݔ�=������9)R
f��+<fKFdnmU+3v3ޠ��E)��	*�W�2� ��fZ�sa`�2��j���!�ȅ$�)�bi-�͠�7ac&K�'̝��ݔ��n�l8R��]����Ҳ�6�n+��k�Ye���p�n��X[���K;e��n��Kz�%-��i��������4[���מo�b�b�@dX6�XO*x�K�}��Y�{;��xyy��,}�C�J��i/n쥾��9�x�et��ޖw��9�+���U*R�{v��+��G�2�p���A"]�C�L��7a����*�#ۻ)w�����<��>ʡgH\��ƪ�$���Iz�<�⬍� � ��%E�����!aKJ����̕y�+D{ۯI��v7r�HE(�P�Z�3"���َ��t�e)=��T�1D:����*%�������i}1�<T�痝�=��w'7�̴���H�D1UFH䖼{2�2U�d�[���,=�������)P����̕̕{wm.�ί>�6�n��<���l��8���� �Nh��J��F���e��v�dktrXj[F7&{=���'�}�KݎL���e_�}yi�iNHDL�]�n��7a��2U�d�X�u�!K��x��Xf�X���*�2R�����|���E)ȩ�J��O�̋�̉o�fZ�q{��W�s�*er��c2HE(�RK�/n�&R̼�����E��C]�J�����6É�-�M�u7l��9��B�$�e���AD�\�e�`W@�l�BL<J[�n�����'>d�~<�IR����&^fia���p���VfJ[~ݤ���������k�fR��J[~ݥ�ٕ��>X�L�*(9NZ��-ݴ���K݅�ɹ>f������0ҝ
$"&e-�n�$�ZZ��I��+�씱��~�_�    ��[Am   &��m��	s�����  H����+f�� �p ��[@ m��v�m�۶�Ɣ��������LL�F9I�-P�����tݞ�:R���6Ա��J�s6��([�f�sg���:KV��W-%��Fn�)i���lK�ic�L;~W�{eެ�U�(��O<�φ��$�';�����*��l����Z-�g8�V���v�v�[��.��.����.^׽�9�e�����_�n�]�&K��@�ٛK���Y�PB��3w쟙3&T���l;c:��	{�!TTq��fD!Vw��_1|d��{���;�H�SR��R�No8��wR�{��o� ����<�i*]�PѱPULLݘ�s3.���T�ʯ���g1�w�~��>��������q�8���� 壄�]�1���ܻL	F�q���kvyА��J�LL7��y�)o��K݆��<�ԢQG�O�̵�$��$!C34��L�U"r���۰�y���:ǖ�����D̥���,3v�2U�d��=��PB%�3Ra�����O�쌋qr�}������$�P��T�\V�c������׹��7a�^f̓318�J�|��kU�fnRh��֍&�:b&��0�R��1##$��*(��T��fD����A��޿d�"�&]D:�$�)��Kosk��7��ٴ�3%�2B�1o��%.L�L��{��~ɴ2_��[����e�`j�zp�^�Z�ۮ%�2�AݼF6�I�\���):��p�6b��� ԬH8�0�c,1%�b$؞/�u΋��a�b�x�޻:�v<"nX�u���D�-��K-�h�<D��5��3-�����e�%�Z`��拢RN΍
X�!`ؖa�͋�I%&"�g�	�8 Xi��&BM!�JNh�yޢ��%<y��ӊ�\xk$�.��
^�����.��.ܼ��2e	&�S��OA�Dd=ঔ:O:_�����|G���s�Ø. _�������	�.,�wo�t�..��7�ڥN�(����)JO|�~�����}��)��>��'.�($e�=��qNH)D!~����z}�����eo|3��sx=�R�{��È��	�{��J>��_o�p�)<�<������漣(���w�[-H��\ 7V�Z�M���5�5M����B]M��#J㳓��^�R����߸=JR#�{���'���~�H>}��8�)I���������N���ӜAĹ�7j�1��JO;�=��)߾�Àґſnm�t��s���֤�H�W$%L�'%(|�<�������)Nb��w��pz��2e�5���)d$[��f����U�k�9������)J_w��p{��;�_}�R���GkpRU��#:D�
hS��=�;�$�0~F�;3ٲ5T�$%R��K��%�������tU d����l�3�pW�<�j=�Gw��YT���f�^�t r��M��Z��	D"3T��B�,�����s���r�{��#T'�kﳊR��w�{��J�}���YrR���Ͽ8=JR�fk럪�:@��9���q{��k���=��y�iJO��߸=H!Kv�]�9�I�[��_j5(�a%�5�o�J7!��}��)��Ͼ��Ԇ�7������JRw�{�%)M}���t��o4kz�@�4�w��pz��>�\R�����JPz{�{�yÂ_��@d��^��_�I���N���ӜA�����������I�����ԥ�ߟ�┥'���������OT�S�%�y����    [Am    ��	4�v�RK�$	�  �m�ø[@�a� (N��}-� -��q��6�m  9nl�a5���˳�����!�p�#L:���u�u�6�R�%�J�.�2������^VMt	�w�u�j&K]vA�e�Ұl��؍"��:UrQv�{�����oE��I;9�O%|�j�
ŵ˕U���V��H�h�c,�"�rM��M�:������ѫ����򔼓 ���=��|� ;�����)JRu�����R��﷥�9���f�d�QQED����D4$^���8��JW�^��\�)O>�\R�����@K�2�j��"�EN��q��&$����R��}��K�2O;�}���~�ÊR���x{��y��:��淾P4��}��)\��<�=������=��)?Ds-I�����R���Y�?�Ѭ�F�oY��R�����JP�)>���R�������X́�gt�L�`M�v��31%�a�홲�[52����Qҷ\�6� �\6���7��dtK��W�'N��/9-S�~���(�~�^�������┥'����R����=�;�F�[�޶qJR��>��Q���H��\[�_���}���qJ}��?5��c�eԥ)��Ê~ �)I�����h�ռ�w���{��;�����)J7����!��N�����S�$�ߺ�PRuJy�k���֭Xmݼ��#K��'����$�\��~���=������� �9��_���Z�	rR����$>�j��]��>�s��͵|�4�>��~��)Jw���┥'�����O,�O������*�j��n���i�M͛�D^M��޹�m�E��I�J�l�B0�;-����5��~�����	��}��qJR����py)\��fZ��.&q{W�Q���8���R������!����&�)>�??0y�2S����R����~��ԞC�������Z4f�6k7���(d���{��S�=����v�g5�y��z*v���=}�_pz��>̚_8��8��h<��F�l$��]^/R����ߟ��������R���V?>����(N��OtnMi��9���Mk]�5A
#�R��q4������)O��\h
C��<�7�'q�d�Aܾ����4�'G�~� m�D�V�-�Κt�uh���R�r�3g��16��s�I�+�6W�Ԇ�%>���qJR��3�qy)J{��┦�����R���V��>jՆ��3{��)I�y�<�y�)��ǯ~�G�rz��{���t)R��'~�Ϯ)��`4���_e�����Y�f�\��z��?>����)J��߸R������)JP��y�44�<���ϫ�-�°��r[�}�k������JS�~����R�0�nO�Ϲ��uPpV_�??:8�)E>�b�"��G)�I$��ӜA�-͚_8�JO;�=�䆣%=��xqJR���9��%������U@WU2�j���c)6\˜�I[�:��&Ko4�*�Ŷo�U����*t�"���s���Şy�r����߾��iJN��߸=JR�{�K��ĸ[���Ԣ턖�����)J}��p�u.KAI��s�R������)JRy�{�du'�.Jy��g�ݫy�[��HQI���ߜ�)��߹ˊS� ��<Ͼ��)��}ÊR4����p��ek7����|�)O��\R������q?/üR������;_|D��>�5���`G��� u-2��n�)JRy�{��JS�=���)>��~�j�R��߷��)JN�>���   hh�  ���`��lБ���I  @l	ж�v�m� 8`v� m� �-�l M���b�Kt�)h9W�fR&�i=�����](p JZGW3X��x�0���G	��sh�k5Ye(�������2B.�e8�Ge V��i�%x����]QO�xy�;9����rI��ʡgH\��V��: 2�T&�-l\�������)�6󫫯U�(d?��R���}�)JR}�����R��߷��)JO;�}��)wW~{��S�Qԥ)UTW� �qo�6���T�ZB�����(J����JR��2��9�]��E��S�����ԥ)��o�R��������?9�r��~~p┥'�}���R���!���P:ADu�.p8���,�S��	.{��R�������P}+������ K�ź��F�l7��s���R��߾�ǒS�4?}�pz��;���qJV����py)O�;�;�����	�5��[:k*�S4Nh���Ռ/1f+���	p�"5��{���B֗y�[��JR}�����R��߷��������qy)J{����_`{x֢�
q���-s�8��[�4�)��zY��a�8.�Ǩ��R���`�C��L��Ϻ:R�������#Jy�k���V�Vw�����&I����<���O���R��;�7'���~pz��P��~s���qw<�f�	UTD����ώ%A��������j����θ=JR��~o��}u�>>��`�jN��y�;y�o9>�}��pe��D�3�R�����R�߿o��ԆI��py)J{���@R��}��Ha��d]M֙�9��`��`0�-e�V
!�G�$�]�|�!����;�Q�o|�������'����R���}��
R����R�ߘ�6�S�GP��\,��5��;�����)JP�~y���@K��4�.p9�[��j5(�a%�޹���)J}��p┥'�{���0�}����0G^� nS�s}\R��-ט�,�s��cXQ*����(%�s���8=�P?�~o�������{�/%)C�~��W�&�\/hfq�E&�9RZ�P)��o�R�~*�����=JR�{��8�)I������R��=���YT,��tU�Z-�`Uġ�t�o	�bP�f���Rvrs��mӼ-�����R���=���S�{�)@�}�׿pz��O�~���i_g���!"*���][\�� 踷7zq=�2R�����'U#J}���┥'�����(�+�=��Z��7�ލ�ֵ��R�&I�{��c�Js����������3�py)J{�e�K�� ��ǖin��s)�K�w��~"Yr����\F������JR���8�4�N�.Ɨl� P��Z�9�~��)J��6�S��wR���qg����H~�{��R�������W8�.���ޗ� �qw���S���I'H�۲�M: )2��󎚪����f�s.� g��R]}�Ԣ턖���k�	($ǐ�~~tqJR�����R�������)���y���ʄ�;������nռѭ�g�)?>�߸=G?3X��ߛ���)Iי��<��=��xp�2R������ѕktk7���)����. �������{��)L��xp�$�����Jϫ^�:�k0۽�ow���&"F���#���}���ԆJw���)JR_����Cԥ�B�}��ˊR��n3�?I	UTD��5Μ�qnnڵ)J?DR�IO���Ӄ�)�~~��.<�Ɉ
O{�=��)������.I_�:!�e����?W�k�oO7�q�ը�XZ�Ѭ��^,DZ?Z�΂bd�Ɏa�#2��8j����7�n�ag`DDV�lI�(����FFE����j0cY��������Ѡ�6Ju�.�ּ�>tw��	˴��8Q7Ĥ�a`�'��s#�8�{BdHnFքͱ�9QubU�Dk5�\ǽ1��l$1����5�)��0B$�4�Y���gK��i�����0A$�����Di�U	$��p;I�A��"c��yӮ����I��ЮզR�*���i����4��';U�UG]+O��zs��wa�f��Ө9{!ո<��y ���YP�Q�rF��5����������\�7*��%�s�� �_��f�St7$                  ������ �      m�                �z   	mp6�     l@ �      ^ݜ�u�    �        M� A��   p         x   �       :@  p�[p -�    �8����g 2 R���� )@A������V�p  �m           � �  ��  ���{:L�c�   �`     z�        ����n�k�X#��<�)Ul*�����Hڠ$�,t�˒�U%���D��v&\�  �r�b��#o��{�A�i���6�5�\mkN\�R���5^;M�5/0�f��q)"Q��L�ր9T�1nƤcCi`k6��b1�
.� �i���[6 �l�MsV�XVW�g��{���60��A��� m[�Jj3((���E�@ �� �p
�����:�f4��Y�������<��u�v*�r@i[�����\E4����b� %��e��m�cL��=��-��ﮀ"
�R4CM�j�F�]��t�fbvMb��u�Dٍ3�K�Ңna�<nWdn�\��-w� �5�&�i���ɨ&�GM1�w6L���t.�Ys��mW.�5���5���R7b�T�i�l:���� �ن��%:ǲ��-��x7z���pN�I �ʒ)@)�v���©_-6�8&�5!Zn5�l ������i�Md��qo��e�\�KJ3RVݙ�q��#\6�^=r�R~��e��|�ԵTz���߽+��>�K�1���|5�?7��jІ���^"�b	��`q>�__ǂq� �/j�j *mW�w�u����{����{� �p���   `���n� �i6 $�t  	 ^�	��0g6�R�����l m�����im�` �3�5!L$Ÿ�Q�� ʕ�5�3oQ��K]�,ܖ�ĻR!%����`��dq�MV-�m�$u�6taٸm`�y���`��X��{V�%c,�M� L-�����}�~y�O<���l8�J�JJ�)6\˜�I�]S����"
��q��2��ݜ�ru���S�Q��UUk��s�L�������q`o��Q�p�0��X�a��7P�8�R9;���>�r�nU곒���@r<�]�]�	O�J�G"�3��;�e�^y�?pIO�_z���P���/ՙ)����q.�Z
��Ssj2T~����߾����a ���З�9	�+�����?+�(��	rLʠ/ݽ~�Iv�R�=�@g�-X�f�Lq�"rUGH�Ur9QmR�)wKT�g�z�Y%��S4\��@�o��[N�N�*nI}nnڰ|����fZ�7��������d��V
�y�s`?u���б_>�7��<I0Z=Cr����E���{�`w�ט��/�9�p�rwuG���DDA)EԽ��ﾥ@��v��}P���vՁ�^���ʣd�S�Qԥ&&f��s�8��?f ���;��U��Y��V�ǖin��q9P�:�=ΚTz3^����{���n��9�`�E.��k�N�m��rsGU������(�+�؂f^����B����;m���U�޷��g�^z9�p��:���qv��^�QRe���U76�����T��y���,���V3MQ��J&
RK��fU���w��G��6�e�	���֏�]�G� ��� 
��J���u�9�32�C�Oӣ�����Q�&A�Uf��~��z���77i�<�>��E9���0s@U��������|�fuY������O�>����|����@�$R��_/"��bY���Ŗ�ni:�LF�l��
X��׽׺�ٔDD�z�׀�ޥ@��o]���K�ή1��v�{6GT�u)JUU -|v�ݧL�wu*r;��Y���$��,�(�C��
��{wm\M��n�33-d���+���*IE����}���7�ڥN�DTr�����	.=��u@3nwR���ή��f��	$O����ء���@ww�ﳖ�ξ����jQ�a%�]��>��@~�O�&o������}J�|��ͩ�����l�ȭ��[T�gKFZ�)���L�Q�f�����WCw���+�g��7��X��t�ɕrw7;�P��5����
��_@�6+��%��n���J�I�go]��$����C'!*�����`{��Vj�S3=z���G�"�HG}�\]�khh�T�(��%(���$�wu*������ڴ�\=�f>X#�>̑�9JS��@B���x�,��T �F�)7�{-XpԿs�@�����o��$�@  ��h   ��	4����\ Hch� @x6�;� V5m�� 2�m ���q���l�� q��]t�����u�֢$ֶ�&y5��t�]��m��v5[�d&�i0[�<U��ᑱL0Lk�f��a���ܼ�ѼHFFs�.��>6խ���b�w4����zV��"
��*�W.P)�'@&\�z$�@�k�e�&�VuΤ��,����'��r�R~����7��6�+1���ե��s{���T����TVz7^�d36�����tԨ)�AykڍJ>����]�������޻?MN�(dϩ��}m@ǲ;����U�L��2��Fq��u��n��;�F��FV�d�v|�ho3�D'e
�f�wu*����fm*�������z���פ��E(����� �D�&�v2���;V6����`�۲N���֯�C'!*��6?�1��{:�\��v���7{�P�s��&QJQqO`���Ui���J�L�'oz����@}�L��.s��&|�۲:� ����)��=�~�	_6�,�#��9��r��`f{mY�g�bޑF���
����J����c�*�0̟���� �`���R�H"*9QX#�Vc�?q����,o�� ��qq���EUT̋K�홲�[52����:l�l�]M�C��Yr�0݈�Kf�GD�wE��޻˶���,ׯ0ģ����G4@�-���;�j�F�'R+o�7��Ķ�ĢM�z����j�B�{��]�K}�R`H�M�;�>��Wi�q%�1�Iw:����ߝ�����M��E���\\�z�0�K�"+�j�mZ�fL&L��Gs�8-��T}�޻fm��`���"�҉Uվ��ޥH�Ivq�V0{w�=8o�t��Y�Ϗ�5�U��Ì�d)�e Ssf�Ӊɠ�|��K�8�1����+m��#�N���
:��Hu������͵`{�L,�{-Xx��"��9N'*'z۽J�̚j3)͞(�Υ@��������9��q�{��J� ��E`�{m�)>G}��zN���w�^Z��R��U-���8�����V����uW���W�/�%)ᘂ�N���>�������s�2���9�w��:��N�V�7�36Ս7��X_o�~����>~��j�
���r �me,��80�Nh��\R�rʲ�].h�,�I���r#����T�Tܒ�fm��}�x��ݥL̙ w����@���s@D\�TX|�٭/�2G];����FOvZ�ˉ	%�0�`~�BDU:Q*���7޻��r=�?f�f�[�Eb�م��>̡� ��H��QZ�I#���b��U.��d�A�L�276���,�(�C��r�Rut��V ��:Pblm*�ݽ�[���H� �d兑a�q�$�ͧQ��˼\@pI�{՟o{�   ��   Z �h�� @����	 m�8'��!���mpm� �h4m�n� ���e����ˮ�WE�`��ц���B�c�J�N.�1l���O���2м�`�6s�]X.���%�Kp�&���/N֍�SA�q�\�;eH+];nC٣���ߺ�_�ڿ�9ӽ�I%UI%2�5��d]M֕ҪI�����5&'c`۴u2��$�S�����7|��N�DR�E`g�|P��ݥ@w�z���TC�h,\��`�uH�z���wR��̹�I� _l��`n��*=��	2d�k�K�D�K��x�T�%�HI}�G�����}J�7�������Vsy��5@H�Mɛ���2vL�w�P�<P��*fI��R��M*3���|�'_4@�҉�T{'J ��eP�޻ݽMA����MeP��.]�+eh� ݆�zp�l���u�ˋ�8Ģ-��9!�lm�����)DԞ�C�3Ԩ�o]��ޥT�gޘXa�e9JD�:��7���Z;d��4��@4��^I�f$���`{6x���ͥI2��yf�F���
��?$���������qG3$�S2I(�ުT��}w�a�����*t�"�r+���zat�ܿnҠ;;z�>fff�n��T�-^^�QRe���*Uـ}��,��=w`>f��=���X��c�d������%�kYn�tӠ�e5L�^+t��y6,�u�]P��c�C�󬜓R�R����JT��t����-#3z�76tM�[�����w~���@!SrN�1�+mZ_�m�XS�ٽR�{�n��A����R*�����/ћ�h�;�n�f�ҤJu���D�߲�ʪ��jQH2���� �MPSO�d��u�	Y�?Y���m�,��,4H�il4�~Ӵ{,�ؖ�'q��b���5Ǯ�)�}��A��[܉'��F$�Fe�!z�����Cf�4��;;��b�l�3F��L�������ght���
>�6�ׅ��a`XY�,�]9�2L��p��,����xs]�0^$`CW�M!��p[$�lM�/�A����a���7�$f��I��4Fi�7�C$t�ť&;��ic��w����}ۢm����N��\_C��������<M*��	�ŗ�р�Cg�D�yy�]��;���&vI߫!���n��*=��:eD"a�JQ7%��Y�|��� ��>Ｌ��T�_��nmq@y�;�yy�K��&��H<�gO]�J��:X���W@ϷvBI*�H��G$�G�RWI��\��L|ӽ�I���o+�^�t3˂R����$�r>�]�n��q9P�;�m���լl�٢��ϻK�2d�2_��y
�¾��������)S��X�ެ-[b�۴��޻�;�S$��N���0�~|���4����T+�%!��닀^����fݫ���|�9���GQ����T�/�C��w�`n��*g�t��6�8i0�K4��!��'�����y��ƨ	��'z��j��G�����r?q���׮,�=y��9�������ʺ�W%s��ڮr�PͷM�\%�~1nݘ��ۅ��I�����Ԟ���'^hDA�Lī�g���*�ݽ{�ުT{ptʈD��nF�;����9��6&Oo������Ł�����/� UG�g��8�u)�U�+ϻ�3;�P2I`���m��yf�F���
���ݵ`{�M,��n��9��^`�$�"����=��
�M�ٖ���z��}��9W���h� c#�"�t��מy�ﾾ��@   ��-���   � !���M�����  @l��[@`�m� ��;m� �� �ݶ &���=u�V�P0��3�����v�����hk�^��5��՗35����)�F�5����R�x�4
������1�j@Hp���/{ށk���\��$S8%}��;�r<�z��l��-Cl)e,��.o/8�d�y8O7d���˃Lg��H�wttK��E�Kݘ���T{�������}���X�<���`�4��55��]�
��(3;�P�:Pk$��Kvz�z����.p�[{��ƨ�7$�����T{'F��:�nҠ��v��`V�kyH�*rTV#�p�ޘ^�/{��~�밈x��@���*!
R��{>?u* I�����7{�M0���v ��.skٲIURE G#�����iyҪI���7"Ú;�3:u,�4��ٚ�WC�AGR�(uQx�{w�{۶����d��c�ݥ@{[ĩw�\޷o{먯<�����U�R���� b�����?���k�g/3�g���=r▿^^%�D �BK�*a)��"^bUS���נ33iQ�d��}�]�=��ŉ(z�i�R��MX*.m`}fd�f߾�&���}w`fl����=�@yfs�F���N�Eh-�ۛ�@��L�I2��������(w��iP#}��5�C�����h��\q.���6��Y��.�n(�j��@� �h[VXl��>�u*,�f��nҦd���o]����sB�ZI��Lz3^���=;��ٛ�l�|�s�w}T�I!�/�K��a��?UD�*b�efZ���*�gw�����O���I&�I�2J+v�mZ
{��v�}����"Tu3*��4?{��l���Tz3^�fdΫ�<�H�uS��	'z��j�3g�5�{v� w�z�f�LÑ��)u��^�tl�ˇ%�1����ي�UJqJϸv�g�$ؖ��Fym�����-�����~����!7��}J�p-_?�49r�)VT���y�J��UUC��0?qdDu��F'��Y�~��{Ư��`*�E*jj,���}��w}�%풲�]�<͖��6�y\j��JUU�"9��Ȉ���/�e�\�>��6fi�4�@t �v��:��,���sB"��f%P��z�ɾa�h��T��}y�5�oM*��Ϥ��E(u��)�r-�N$�u٩�[-t�i��f�X�U-����1;/`fwR�;ݽv&��T�K䐙$�<�5����8�*4JTVϢ9
�n��RogZq��q|�%�s�\\L=�-��uS��#��5���@��z<���T��]��{������\K��.?�ⷞ��Ԩ�w��t�3����_��3���r���<���V9�K�.�����}J�]��zٙ��2Q���Ͼ�  �m�   �lU�[�t�K�	!�(  ��$ ��6؃���� 6��:m��[�UUb�E��h$�ɒ��!#�3Mb��C�T�p��Y��:�%�Af�m�4�-���{�^���0���ktX��ieM��PbKp-�9�[്���t�A��ճ�_��=�����:w�
�u`���;6�g.b�2�����Y]����L�
4��(mH�u�s��Dr1өQj~���@�۴�ލ�fd�@{ٴ�1������u L�D��ڰ=�ԫ�b�R��7��T���ԩ#���I$�	�4" �i���@w�u��fҡ�;�n��{v����@Z"�D�J%]�����L��2K�37WߞTߟ}�v�wR���⬟��]�t=����"Pꢰ��۽vL�/gu*��@O��j�?}����k*�tR�m[Mf� �su���i�e�&9�`�5�e��c��Ո���3�� ;Ѻ���J�33~!4s���a y�	�"��
������g���:SԖ8 �/��X>+��q`??{0�u�ZH�����%�R���{��J�������/��9#~�q`~����F�5_)D�J�
b&%P���`���Tz7^���ɾas�/V�S��}�����j��
�I;`{7�T;���z�ݥ@on�ߝ�]��@�$R��[:e�M��:�M�e�lsH��(ʃ�Jw��'�Y9�yo�[4�$�(���	S�
Ϸr0�o0��T{AptʈD���^�^��?g9�Gk��Y�n�\Xu>�j�8`}��%F�M�E|@,�������1�7ČL��N$�6F2L�@A0@�2F-�bLAX���@C3$A%��	,�HG �hG��y��{9�#�l������z=ϊ�;z�R5�4��T�Ĉ)�J�*w�{ٶ��<�ұ��{-X/s����{����	�"��
����N��@3&M~ݥH<�ѽv������[�~j�
�\ �M��he�m%knM�b�4�Ͳ�Q�1�7���/z]E*����fwR�p~���f�*e�.�����fs�5H�:���{d�>vJk����H�N��rե�qM��۷�T�U*Iއ��T�mq`/gu*{7����u��US'!%Ea�%�qqr�~�^���y��Y��u�qC�
T$�_�ē\�S{[]�`nxȪ�)҉C�
��wR�>I���f]�����;�V���=�^ɲSrH���t㧐���UU�D~&�흤�[��ZF%��f�w[��� ��R*�uQwϴ�����fnڰ7�L,߳-X��إ:�
R��&�+ޤ�P��ԊL�ݽ:V;�~ͻ]����&�1�y��M��T��͝(��,V�tu2J��{n��n�R�Fh/,{G)��U��/m� �^ڰF�o]��f��#3��t�N�-��z�QIʩQ�73z��s�K3ut�����J�c�//���i�@_� �����C���	� ����Q��r7��`��u�j&��ȎX�7�Ր$�n���JF^/��B�.��p���n�������u�����5��EK���dDkXM�3 ��'�S@?�V�yE�`C6�a$�H$`��Xd$�$΁�l6��߹�(�����I�	�%�Bd�����B�5�d�&
n�I�׽yݣVk+(�V���h̍Q�j�8Z5��7f�e樧"�.���#�aWAJ>)I��?�{�?{��M-                    m           8                     -��n�    �6��m�       [��%�Rv  �          �m� ���               N�)Cm�   `H  i1      �\�A��m�J  d �� 2 R��հd   ���            ��     ���ֵ��  ��    8           mw-�6�U�B46�qE��_��]ѝ��y�!\��	��S��;�s�W43�hZ�ʭ���5K��3g�W���l�]�JZD6�g$YrM���!�;��Ub�X����bX�6�";�/�n�G�j��%���/�C;\b6�U7���,�U!!X�l5�>y��ݾ�oVڪ5� lCpIf��Wf(LZ�v��غ��e�-p����DrK��6�s��Hl�Y� �e���[��:��(a�2��`���X���(wX`
UU���j�\�m�uԳ.�8���pE����I�k�W\ L�R�kQ�3]33��nP�b�ZM��4ѵ��.�8�el�ϧ����{='�_��Z� ����[F:Yn�h��`&C�	vŒ�Mui5*�k1.�9hg����H�f(gh�^(FWr�R����^�촴�GlR�w��R�\J����PѮ�����8�5	[0le�an���Y@�R�~{��iqxSs�h������36�3�9n嫣tЀ�bΦ����ξ{�]�h�H�ј�� F���粟�:��9k��YM�x��"`+��ЇJ����4o�����󻻽�/ϖP    [Am    ��	4�����8  �����-�]�6����ж� ��Aƻm��  s]#�}�=�Z��]��HM��a:t��)���ue���u�5��b�f��vKyq]��l�н���l���Af�K|^�wF]�\f٥�ZR�gJڲ�v#,�m�P�m�j��|������z@����[��4�6*)T�]���B^XgT˵��bl�h������/h�ԩ w�4�/۴�$���t��n��:��䴓1*�����d�L�dc�iP��[ێ��֫�̙!��ۡUD�*b�%e�@=~������rmQ�z���j�w��Ƽ�ȩML0��E��Ȉ����~��f'�֨�������7�0�"S)T�*��;�w~K�t� >�w�~}���'ߟ_HaA��k+���s.sm&l\����^��%+i�lrU��r�e����AJ���d��.��k:��o3 �u�\g#��e�"���rQ��n.��n�>��6&� <8X�24P�X�u�k#d�&lR�d�̕�>^$֗���v�z��d��>Y���%(
�NQRr����V�z��ӦI�vt�@�ͥN�{x���&�UIހ���V��l���3mZ
O73~�l�g�R�UD�$Ī
��� ���ݥ@۽V�z�m�}���� �j��u�9+m݆�zp�g-�.��L�fW`%on;l-���1�L�����`?7��>�w�BF�L/�����mk�AGR�t��V���=	o�{��w�q`b�?j��A)Mʨ���fm�:��On]���ʹ�������'�{�������}�־��n����17H"�\�k���&O��q@{w�P��\[��^��V��99(�Q7SWF�븶��3{����kz�����^Y7d$��	�5��[:i�m���Nh��Vy.4�u�X�ۏ��{V�$m�&J,�������������mi����dXѦ�Õ\#���Rw�}�������%�k~��V������\?hM�_�J�U����w=�4P�����:7z���T{ptʈD��c�xL�=�J�����z� �fLڒ���5� X}��9J��UEh�;�Wٛ�d;�l�
�=����$��}�L�31'8�n�n���ҺUI	�X�����R"8�SJ��o/��!�M�H� ������?���3�ۉ��T����# c~"o�j]J��o�a���$#۵J�[۽v�z��?@���Uj�K�@�3mXp�������3m[l�d��_,�cw�J���T�Ü᛺� �u�X����;sݧ�`f�4�h�%�:����۽J��l�@^f��7�{��u�z�$���K���Ͽ]w�   [@[@�`   � ��M�$$ ��NR� Hm��:�.ٍ��,� �  l[v� 8�J��P�p��m�m�-콁�u ��$�Am��Fm`b%h�.4yJ#�J��p����/{���6m,h����^8�3�-6"��1��,�0��R�K���C����y���9���B�X T�@�T��^rI'3�r���8��*�[`���6�/M�Vvk(�b��WQ(9�
�[�h�P�KI3��}<Py�j�7�~}7�fe���Fw}J�n7��ʈD���]�w�R��h��J�߲a`4�ec�A���S��S���]���J��B~��yS��������m�uv�9�{-X�3� ]��X{�2�߻��!ϑP��J���T��(L��m*{w�-��͵h��l���	T۪��bU@(U�s��y<�MLxF̲7��I�P�v�h�5��J����=�Ԩw�z�|�2�]��'�#��h���cw�J���T�Ç����]v �E����v*ww�;��ĥ�`��,�j|"&xR�Q53U��}��/��S�Y�"9:ۨ�;۽v�#Y�4(��%���T�l�@g{��ט4���XRt!����L<)P!�E���J�2K{w����ڰ7����X�sd$����@��-��Ȧ�J�U$�{E�5a5��4@`%�fkmA34�UUR�Sə����`6�+{B�0������}�f�)�R�ܪ�N��v��\\���K�C�n�����V~�oz3�{Z�Q7H���*���z36�#�M���V�̒�Z�^���{��2�L��L���V݁��X�;99(�QqWJ���s�M�dXp����ͻ��{��r3�~�1~����%(
�N'R+73{�8��ԩ=��{^fҠF�7�aǗ�:�.譼V�j��K�X�7&�v��m�6�n(�\���Kթ\g����h �yo��߿y:�Oݶ��Kd޻����xXV��*��'(���7��w�s��R�\�-�q`?7��>m�Xpt!����L<)J.)���T!۽ve�32�7{j�Y��v��+r�9N�UQP۽j��wR��������%�̙'J"��h/P����xs���foҦ$A
a�b��Z��h�;&K��|�n�R�73�$�ٽ2j*�\��Rʨ���VU8#��3���f�PE�#ss���lJf ��[_e�n#�H��qp�מ��w��ŀG������ˍZ��}ffڿ��5�H6���Q�{�}-� >��jW�J���Ԋ��n�����ڳɽ�m���Z�G�1����MTrN�r#�6�,���b7u�<Mc��o�AЬ�[�UUTNQ%E`oպ��&d$�:h[�Ԭ���=�Ԩ�s���;��|����d�    ��[B@   ��u��I� $g@  ��@�̐6�g6�2 R�m�` ڶ�����-�l M�5k�,r������©6 L�b8Ylh���������6Zh݅5r[��G�0𛷻�{�h��Xq�b���,�$4�6�Sh`�\e��n��kh����	tq��o������$���l8�J�|��kU��H�h��8�e��b4��U�Z��ڬP#!����O����{���ͼ���ڰ��u� �#��U����{��z�9�P�~���G�=
��3iU���k�S �2�L�U�'��E���e��{[qpg����a��+X�&�(�REa�qp:e��u�`w^NL��m�Xa����e(���WF�����y�[�wmX�f�6��eȤm�H�9\������T]YY�]�`L�(��ء�'��}�9�5S���R����u"��*n������>t�G1ԍ���Õ\#��*��@�wm\Is���%j�_MNfm*��뱒�L&Ng�3��DD�LĪ	N�>���6��1�u݁��J����L����R�=�t��r9�\�q��w��cH�qa#�XC�q�"H�:�UEaO�w�gwJ�=�(��T���^BtR�m[Mf� ��4ܭw��-]���0K���N%�0�igL�|�9?�fpϾ��3>��ffҠ{���ֱTM�Q���}�օ�ffڵ	�����6�����2P�n������e(���WFr�y��?X����,�b�g�×��А���ե���Bɨ��@뮴�̹��e�LcZ�w�~���Ig��k?H�kZM�Xe�P���[�h*�F�գ��5��I�e����b���u����΄�i�~���Bƫ��R�8qx	�16dĪF���@�4=��,���M`ê&��Q��y�;�۠8$JLE�퐒�m`�\��ڽ�l�H�"8ҧ!��n��bܝ����a�s+=U���A� t
;��$+0C�zxhQ���� O ��@�� ��Mf�᫭��ȧyϿ����Y�S�����n�)@TRq:�X�w]���@{�<P��3�m*�k�|93B�&j� ��j��|��y�<��۽�@�{6�$����@�L����Q�e p�F�G��;�Ym3H��\��"A'�)U6NQ*G�>�&�#fKV����p�Gs�����tX�ԫ�%q�ﾻr>��{g� �}��9I�JIa���zy����m����{�,�LOǳb��)�n���������M;��2s�����E ��C��>�?O���O�,��*��
"�R��>��K��X�n��Wۻ�ߝ�*Mzfl$�������"mL�@s.sn&i.v��HA4���U�1ҫj�&��9L�5j\r���wgP=o0�w]��"�4���Wʘ�PBy�����k�s;���d��Ё뺰;�M>��J�D��V} O]*��![��&d��>��΂L��ƺ�:��_(���~�YK_��F��ݸ?��v�z��p.�Q0�JP�E���>e��>pϻ�T��=���
u�:z�A$)Жɤ�������Nr|�/�~�����I��[@  6ؚ�	4����l Hkh� @x6�;� V5m�� 2�m �6���T�AUU���t1�&
|�:wKsV"Y�6�ea..�-�մ�;�+v{+��h�s6���Y��sm�MʤJ�O"t�œ����K���h��کA���bƹ�M"�զ2�#o���C�N�9�\������SrH�#�ꮵ��i�M͛�N'&��D��D+)<p��U��GUr
9*S�
�~�n�R�nm�����V�;�oM�7��0�"rG�S7d;���V2Ob�^ʎ(svh��v3P�<��(�%LDĪ3g� �f�/���A�ޥP�<���eƭK�\: 33e�}�7��=w�{�,�;�|����DL���v��oR�N�{�<W������v�O��~Z����\�;YK*�\S�-v�&!/,3�b�`bl�O��{��^�DDL߄�Ԩ{'� �f�ɭ�fI$_�߾����u�
%���\����ֹ�� I�!�w��N�}���u�Yi}�`�d*T�+,���XR����6r�Ł�ޚXCެq�(�(I%���u�n�����zݚ����n��N���*��� �͊�6~K��_n���@?{��b9�Pw��f ߫�EUT̎�n�YSu�t���q\��ƭ�X���ڱ�ˋp:��Rұ�3�|�ܞ(}�4{��~L��>��� v��yzNJ.�\Uҫ� [���!����o�>�9aK��楜��L�QP"���hv�R�}dғ-�֦d�37��se��ե�c���Ip�v���4~}��3��7�:PS�7�`fk:�	�b"QN�<[W)��,
��u���q`~�r9�=���U:B�ܲ�V� �� �M,Wqp1�aIY�
�d%2����6�`Z������_�ԍ�y�'��,}�Y g�̢IBE\�����������W����g�a��e��M��3E)� &(�%5���Ł���#䷻w�gG]�x3��Q(r��J��I0��l�S�gu�����s5����	����H~*'�t��~~wҤ߁j���uJk�*��y��֨�r��|Tr�~��>{L�#���P-.�Sdv6��U@�Sq�[��:��LGKj���ۏ�#����Hm�$e�%`,�����o��{���1�Y��r1@>�qi#�7����A$�l���x��T�&dߢhr;��w~����'+a>T�(hwxR�O��RC���n��ޥ@caTLLT�*"VY�B�!{}��|���u�lF"W�o ��d٨Ԫ���UQY�����@�ʹ��}���Y���=�U���,`�)*<��?��[��   ��h   � I�M� ��� Hd� 
T�6�;���� ���6� m�n��.�UUV A�����]�2
�;<�8���4m1�Q������h�ÜJB+��UvL���ny)P��)z�t����ղ���9^JY%-��D��pʴ[����w��{�U@V)@[����n���S��
�-�[�[);-m�0h?�qR�-Jj���*����o�֭1��`o�ZX������-4�!0K�īݳ��}��������k]��Hބz���c����U�|���X��a興���W�����~,�7D;�L�!�"J�$�s���o�>�,����ݖ}�V�Ó0R	������^E�Gߣ��#i��ե�ouᐁ��U(T���T��ە��.�Izh�i��mK�.��ua��g��|j��p�J����������_R�^~�D|���߲0 ��G��Q&��5l5�r��Ϸ��(>7`=�|��r;�{oـG_�p�7���o�ܢUF�T$Uʩn{7�s6՟�?nU^�u�`y{���-{{�èR4ď0�7`��w�Pܝ2��Δ������*�e"�ӨX�L/��Ԃ{:_ {�y�>�e���몜�V�j`qK)eT�G	��ja#Z2h��#�nn�N8���5���ƭK�\:�M�@����L�#9���x�;���H��DUU��f����u�Xݝ(���~2ei����I~w�&+�����/rt�s��%����/ѫG�����뭟��	p\I:�}z�ax����ށ��g�7\9Q�>=0�3ޘX���@�l������*R�*Y�+s/���K��{�;��O��d�R�|���?����@�$R��_/"�˙nF�Ia]R5a4��71�8i�gI$,4l��!Ф��<���`vt�@^��A���?���L:� CLH�����|��r�J�� ��ӕV���y�@gX�&�"�ӨXu��� ׹���C�뷙�>�fb!599(��`ȼ�yG�=�e����)#^�e�܊�9�rs�2�����`��DR"��X{�2�#��r7���i�7��;l�}����ڹVe��٥pR�$kVx�����MoR7qfu�S��KWlJ&k0��F���H��֟b�{�����B��jn�A �7!`�}�J@nd�@v����(���*)N��>��fM.�7=�ޓJ�˚X#�0�lFc3h�Q�U	r�B�����L9�����ҁ�e����9ϳuJj��*S��Iu�۳K۳�����f���g�~����C����2����w��D��PE~����ց'�� S���I�L�8�-4Jh(���'��'{C��H�6�AN�,Өlх�e���/�n;�����,�g*e�h�����F	�	�C� �H���4��ډ��PE�a����F�ѭe�k	�f���B�ķs]i�s_'=�!���5���<%45�񛢭�9�5?]ǳv~����6`��*�                   �         6�                      m���    p� l�      ��i��          �  � �[@N�          �     H �    �  6�X $     )!!��pl  d �� 2 R�����b  km�          -� [@     Bu�uv��ڰ                  �`(�|�i+������w\�y��_�x�GNATr��I���!�^͉��[S��4h�"\�n�.��R�G����x��j���x]]�]zc�Z���+!(N���7^��78֎�H�(�*�m����# ��Ei������L̎I���fΡ�Kˣ5�iV�޾|���}��*��[U]��e��*���e�4�ö[��B�l�2�c�6Մۦ:dT�H?am�ބ!��\6|�Fx�G$�qX�V^4m����B1�Jg �AbU�n�������K;�+��]`9�
[CE&�q)���Pź���h�%M��.�`���������n�Ujk`�@�����ϓ�ϛm��͵ī:�[�-�.k���Dqtķ�м�gA&n�;�mA�h�lۥ�.�jZ!���[+�S6l�5�����[6�jRSq��v��b�&�
�ۣic-,rݶ�M�b�Bf��I�c��U�a���&�β�h�4[�m�[�J�2�Y�����p`Q-�mL�����2�&z�����4���D��K�)�UJ`���w���ت�S�'��*|�lOP$n��:6�
@�����w����{  i�[Am    ZH��6[����  @l�8�����`8�hv� m� �-�l 2C�sr��K���\��R=���X��6VT.��鬰��#UY��u�����ZjM�4�l��ޫbDl������s-���JK`��]�s��^Qpk�s�s�����'';<���ֲ�zi�I�74��l�S��a�ˑsF��Rڣ��%��������Y`n�2�{�y8���4��P=qk�hr��)˨���>�k� ���=Ι`��m��G9�L��%|��f
��������>n�e%����&�v�f��4��ɘ
��(���>n�p~ݩ(̝(32~�����8&Y�'w���9�鄶���n��~��}��?�w�|�� m�)@[���Mj�,�ɺ�m�RgN�z�Md���r�􅓒���Q53��$���]������Is�'ۗ�@3�f�*�R�*�T������X8@0Hb)	$��F �ؐD�A1���H�L�8��0UP>�.�C��~����Ʌ��za`u}��ST��Pr�M��+�n�fN�no]�x=��Uj�R�T��W��޼,�����gb�{����r=#Q�������WF���)'�ט^�,#�z���#$mԌ��rW�6VI-R�m�,H�ke��`�t�SQ�(mH�[0Yvy$@U"*���{����{ria��̻,{��9��1���A#l�UN�wO�ϓ����ۛ�33�����~M��H*#��fz�۲����'�P(VV �%e�5�4��"�#�W���<��O�L��)J������ȈM��`y��`7L�����ϧ.{v�7����J�Ԫ���L���� ��m`=�X��v��=����*��Ä�����I�su��a����W�=�{N�5[i(�4#m8�<����{��U�����HA��@v�oz�{kX�&�"��TW��U��3܎s���֬����05kuq`?��p�����qW����N�v����$��&��kz�{2�>Y�!���P�/A��vz�v�*);���G2Y���S�U������U�w��>��U$�D�fZT�z�,G7vـg�5�|�fM�B'����I%UI��Uv6���(�u6F:�bKi�F���qSHq��댐TJ���&��c����zۛj������'MTJg,����j�ɑ�o0�]Ņ��ޖ�fe�5*�6�仏�w=���gs��X��*g�5�������4��^^"n��oR�/wiP��z���Ɏ�査��|����`���jj7G�v�>zs^�N��޻gwR���f""��!���L�5��D�L_y��k�����  h��   m�MV�n�i. $�h� @r%�H<$ �g6�R��m�` mmm[�۶�ƶ����M����H��Nd�FvЛ0ۢ���bbqn�ΖK����9�"I�]���V���X��,S��m�Η����Eي[�X[EnB9zg�w7Kw+�|��þ�9��s�����|�U@WU3cmL�@s.si>��ٺ]� M2i��ȅ�L��StST��r��;R�r�@�V��ޫ|��TnΔ��w����������I=w�G�5���=���G8��55����I�Mf�?\X��>K���`=z� ���jc�2AQ*��3
�����;g7^oN��smX��ȤQ:j�*v����֯R=�z߾q��]��GvwU�-���|5�Bΐ�r[[Mf� ݆�^�NM3�7����*�<B%��a�t�J��Y<��XM�����/�J���`w����ʼ�S�����7S��͵muAE4444[~���Jb�Nk����L$o���@�������2��{�`{[y�%�u�DMBQ0MIS55vwU��~����&������}���l�5�M�+��R�待<��v���L�tDF�*�ge�-��M2 *�:����ށ��ڰ=����ϻ������媠*��UPck)eTˁ�sE���Մ%�:��Q�L�1u1�^	N�u;�>��R�{+1��yU�����>a;����(��j,����נ;{��:�oZ��{48:b���r�n:Ϩ�ih�w{ѯ˝=|jP�]�J��̵�ߚ���Pə[t߶��Fk�c����&"]LD�*&e�9�&X�C&����`C3,����=��v ���v���USRpDNH��?�g]Łݝ�a�{[i����'ϟ_HaA��k"�n���RI�x.�ܑ	/N�Z��\�V;~�m��`͡-J%T��ͭ�`fzdv������_.|�qm#�5�K$�9J.*�����V�I_�����;>�T�0�׽��%@
�EN��l�f~�P��V(����c�;�{�b�<{�U �(RJ���]ŀwV�K�Wuf"y����7��bh-}���޷��}�T�Z�T'j�U�ܬ�`{��<��7{�ۛj���vJc�I�GK�:�V� ����zq<���8��(� �!(��p($�H��ʝ��z�Yl77w�ۛk�gee� ���Q*�R�*��Ұ��&/�^F�OuX�wU���=�TԜ8���@��ھ�T���V[����x���y��F�M�&��A�LJ�3cu�V\��נ=�s����Ȱ3�A''	�QqWuk ��j�z���]Łݝ�`g�o��   $ ��-    ��	4����l kXHh� A�m�8w �fm�� )m�m m���v��[@ �c羥���ug'k�h�Ӗ��"کn��Gaԩ�ˉ�[6�\U�B�h-r0���k陫6���sntn�l�$���,o�.�v/��t����u���~��{�xs�9�Bt�V���e�[��4�6�MS'4b�F7Yqt&m�V�A-�����b]�#m�+��ٵ�'�9�a0��]Łݝ�`w��V�uj|9T�FӢ�����V�����՘�)�no�-��+8֦U	��UD[�f���ףnf{�z���T,մ"�@t�NT����K�2m�ss{�7�V�{/-�y��J�Ԫ���MM+ �y�u븰;��V��>��}�|����H�n�n�2�e̹ʹ��,#Ʋ�H�J�tfI�G��l04^Y^j�J�3䎺wv{���Ӻ��^g �
�*�mQR�U*+�^�{����:���D��o�*s{�޼�`w��Ƒ�����#�	�S�'	�QqVV���ϼ�o����^�g��ɂ�J��*r;ss{`goR�3c5��n� ��;���i��U��e��u�}�Sj���y�{���=Oު�*UUH��f��V�+E�
]�j���߹ַ�c��tŹ���a��V:�8�L��5Cu�׵����_�ٽ��M,��CdQH��*v��>춯�Ɏv��_��@۫,��U�9	u.�5�S4��h����Ұ<�����zt�k�&�m6Rbc]"�T�6�1��Z�ka��
(<h'f[�;І�/�Q��-�tJ�EGkP</8�`�d�yQGk�޺�Hc�������p$��T�Z�3z�5����A����� 6����{v#�*B�x����J�>v�������M!�1�^]lFK/+Lɚ�t�F����z%��=�TԜ8����6�eM,��z
{��xL�H�����7��eN6��D���U�v���v�{�=�X���?o�)�%UI  �CdqK)eT�G	ɣs
vY4^h�4)��;WZ���_LVA��� �ϼ��^`��r��^�`$���`�%Sq��T��^cQ�ue�!l�U��N�M�����R
�N�rv���ɥ�ܞ꿗�)L�U����29�/�V�C�G����Wl�vO�L�`w7:�.� �2wd�B��y��;���T��r�����=�;�`|ɾ��xޟ��^�q6u<�HI%UI��@[���Mi]%d�u�2qۯN^����Æ��,�ܩ����RG�Xo�����^�r���o�Vk�ki��ߕSRpD�7U��Ou�3܎A�[Vݝj���y�=�TeN6��D�������~��1'-��>��,�բ�')D�V�#��N��S#׏0�i�	��v�{7|��P%:�����=�<P����3^���)��Oy�ν����_��w��޿    ������   -hM�S`		  q��� $����B��1��p �E��� [dA�ݶ ZB��_<r4[����W]I��P��F�Um�,�δ1��k���+��wQ�LB2J�a��;�^�х��[q�V*4�xm\h��2�h-��t�b1��*�n:� +��|7��o'�rNIg$�ӻ�=Sm\���y�+E�J��,H��M��)M�#�(��NdM����AD㢝O�ٓ�g�yY���Fk�8Gow{�{5�s<("^]@��`wguX��U����`��. �f�Ȣ�5S�;q�:���w�L�[�¹Ȅ���,�9���z��:��NT�UBE\�#�77w��d���Vc�����vW��USRpENS����wi�vwU�#�&�Y�7Z� �
:��ePN�]k.צ� ��sJ����q���j�h�Ƹh�3mWQ�|\�V��ֵ�o�מ�s��^,i����')D�/�gZ�G+���
YrfL�bO������Mlf�|�!)[YYʚ+�%X\���c��0f�$���ci�2`H��潁9���Ó0W����<����ε`gӺ�kן}������1$ҥ%4X%�WuX���^eBG��e�������q"���ӑL�n�F�E�f,�����e���ڬͪ�1��x>],��j�z����3�� �:՟&?36��"�P�R�征�7w���������`^F��n�s$��̓^���jN�rF��@�����?f��9pS��O�W_�� :41�w%��DF ׯ1��:d�&�$H�J�SE����T�j�K�Kk؁|�����S��<XJ�Ʀ#�p��D�V�R;�mX[y�w�L�b��W$�y�}����`��o-f��n�\�.������|���d���+H6���fvx�uS4��T���y�W{��6{��Ȉ��b��ڰ7�S^�ɘ	+�IUY����j��(C��V{-������kx�QQƨu#�=��v�Vc���dٹ���7jk�>���(�L��*e��;�mX^��;�m]B[""i��9�~�`�=�ܩ�	J�54�7Z� �[VZ]��#�����ݶ�����5�U�.&�5,�
M˛��}��=�,�t����?vtu�V�Je���i8� ���o�M�`/e{��՘����@0�ң*!�C�J�#�=��uu(���V���:���6�ӫD98NR���]Z��e�`f�y��]�~��`g�1ݷI�f`7�J�c���ꕁ��;�mXp��uY���*"�vڰ:Φ�Ó0W��� �e�`wg�����`=z� ��Ȟq�HwUU@  h��   `5��p	6�`@H΀  ��	 `�m�d ���� 6�`p���ŷm��q=��c��7]%�湎�,�0�bˡq�Yu��\q3��L����ú\g_���-u�4]�U�]X;1��1��p,�Z��h촺���P�i��?Ru�F�R'w��n�����9;�N�*�P��P�gL�i�˶Y���c��Y�/i;AR�ط���|jqҢ��P�G�_ޞ��=��;~���@��u�&�b�dQH�$�&��`춯�:r�Kv]��^�}M���e7*D�R�T��
���xY��3lf��F����E5" �rF��@��u�n߲{�3+��#��ߺ���*2��M���JY }�ZX���i��y��0�[��~~�����,5(�[��lԍ̹̤ѱ�.��L�3K���x�c�lST����m�&��;�j����>]n}�A�i���%|����i*�Xׯ3��#�|UWA��NY{���r�<�\�ތנ=�>�0� �x!�n���tY�#�wv����&����k ��y�u�g�:TTqӪ��g��W��u��˭́�abbf$�&�(�;�֬���]��-͐Z߶��>�����Y�.Kkeh� .R
��ű�X�i��.f[��t�������t�ebC�̽�úw��S�gtP�1[�di!���{����7S����1>��Xb�OZ�;���-i�ɤM$��G$���^�ް�IX��\\R���yO��63/2I�k��2�Ͻ�h{ͼ�p��V��|��&��>Z�y�����zp29�ו��	N�K9SE!L�*TҰ7�7�GW[�}[��������f�I%UI A6�n�tӠ�e.�o/l�na4��䩆`�b�"Zʕ\93%qL�k0��64�e����[�nn��}�YƷ�ES�j�I��;���q!�[V��� {:Ձ��[J���T��}�$��uհ����ǹ�%�O��l�� 7�j6�D�JUʒ;��w�#{��v�{��hC�~���IG�������-����#����@�B:��=�j���N걤�-��?���>|��@��n�YSM�2�6RX�e�fe�V
4gV�ZX䳥A2��lҴ�ST���VDi;���3�� �u�{Ԗ�rp��6uk �r!�[W)��������wU��ކ��M$�i*iṂ^��rk�O����wV��U�Ó0W�SY�=�j�}��`oӺ�=�:���w��k�*���J�;ے��6?�1���z�p��w�!�!	 I�L��CD�ㄑLL[ۍ�ևZ�.&��V��54P��Xd�o!!����M����n����A��z�8@�Q�;z@�T6ȝ�@j)�
*�1,5�`���Zx��|X����!B�l�J$�b2��sM��2�j�m��{���[�)�qy�p��k�!����|����e�1K�7V��
*&7�\�W���&�h                    ��       ��?�=                     �l�    �m�	 �`$       R��5���            m� ��               �       	�� Hm�� A�  ӏA���@A��6�2 R���� )@A����� Z� d  մ         ��� �    � ��e�+�ƺ�                  �`)��ش�h�1�f����;|��u�����(����<�j���3��#KWO�\��]E f̢W)H�#U��:�6օ��`�8k�U�6́��:K��n��}��$CH�B��$	b��(�mƹ+v�9��M�0K����9��	��gJ��QR��ll5$����w��E1Jp�$�GUU\�b���-R�&��h`U)����0�`�F�m��@�)�����%�4[�([�Ӳ��w{A��&�V�ۊ�1*�x��v�\�l1��)�-��!��������#j]�lssF�%�	�����ڍ���YMtT]VCA���b�$�6-[j%\�@�sW_�=���	|��M�f��ۛ�1T��h�SS�.İ�r]Gܥ��6T�j�J�I+rV��&3��D65�c�Z�'�\S��l �ʺhM���]V4�6�C!��n�v���um�_;b�5Lv��tMJS5��g�y;�d�0�[�ZX`�#e�5�n�[6��`vi�UF�\�ַ%7���}=�|wç�<�{�{l��^���N��çrBA8��.y�����k�7�����.��Cv!�+�C��Q�1OG�@S�t��M� �>:����{����{  $ ���   j�$�m��I6 $�h� @x6�<$Xն�  �(u� �[A�k���-�l ��,m�'׳�b$�ɷV��TmSMRS����֦X�����5AkL�s&؀kRF�mz���t��i&l$AVl���Ӻ=�i�̥<(	�X�(o7z�[�]���+|ݱD8z����]u����y��gH\���eh�
]�c��w������̮��0 �IE �lHLmiG��u��~|>�5_ҍt�`�-���X���~F�j�N)�\�#�Fnn���R=ھ�l7՘���^�`b�=�TԈ&HG5���V�wUZ������� �7J���eQ����[�&};� �m��Ԇ�ڴ��u%��')M���Z�gZ�?�������{e�n ����Iϝ��骛`��k-�YK*�S4Nh��J�l��B�(��v�?��wY��x�D��"�U/�~���^ԵgR}���qpa���`f���|�"eU9;�gZ�9��ڰgZ�5��D�L\��+x�~䄧#|�$�����wԍ��>��o��`e�`}��j��ʂI�T���)������m� �u���7�a�3��N)�\�Q�ׯ0}�j��^�~��	>����E(u�t]M֮e�m�ЬɬYx�YH��D����t6,��j�����W)�z���R�"�k�y�L��ۥFTM��(�J��[�f;�fvvՄ�^`��3=�rL�u$�zN����n�`�~WI�^aq��:, �I� x,�p�`�LM��=u�s�hx��+� �[zՁ�}^�`yg��T ۪�����Z�_��;��3�V Řc���� �N�rw�&�6�]�z"#��y�5.��V��� k[��%:.譼V�l�K�շJ��ҫ]m�-aaJ8�
�[�h���4��o���kSh#z�� ����֡LLL��\�˥�>ε~�%i�H�����{�.@��fJ�8�Nʕ��v���Ԩ�du=��נ5n=�TԈB�R�ށ�͵`oո�:�s^{��|�H**b���P��� �TLC��A5ľ�׻�Iw꛽���TeD�(n(����C�V�=�`o^��u�Y'�w���᪛`��k.�tӪ�Z8Nh�ܡu�+�Լp�V���fTM�uK�z��V�#f�� ޿�a�=wq6��/U�՞w�P�n�2S������UF�6Ս����q%bI�>�c���3v�)r��*D̪��u�X��V{��9�0�ߜ��}�{3 �	�(|��SU+�U3Q`?�uX��U��u�]�w�����:T����rWn>�?���5��޻��J��F��e��dƿ��w�   ��   Z �H�l)%�@�N  	e����-�m����� �h8�fl�� �h˻Z�}��_����#h��Dp�7K���锛&e�&w����[p��J��]����k��p�Z�MSmv+jRX�2��[K��.G�u��v��D��6��:\������x����V���[�-��Ȧ����Hv�Fń��LD�j����{�m��$�N)+�*=f{?w�}��,��_�#����j�p�{�2��"�R�UV`u���#&$~u-X��X�7{ߒM��TeD6�2)$����z�Fk���ގ�=�Ԩ	�Ė�rp��L\\Mկ�ݝj�׭��[��B�����5|�����"�M+}���sw���=�ڰ>�wU�u�����i"���y�+E�˘�����]a��٩�mD)��1�̝������r��S_|�wb3�����ڰ��w~�Ь�Ox*�RSUNTV����! v��
:;{����>}טz�t7Z�10�D̕�Yt� �e�bK^��z9��=2�W��X��]�/�f3$�N)+�$v~�y�w��X���+n�ܽV�u7)H�(�G����~��웯��~����6�w� _fl���A���]�M: )	su�輆v�.�y�T�X������
���*�)$���f;�1�׭�[��\��KD98NR�����{2;��3/B�z{�ɗ�+w�Ձ�^�b^�c�J�uQ��Gzٵ��uE�y��\���K��TUM�HH�� �I���؜fT�&񰟣q���z0��揕GUN�z��j��������v��`�N�C�52�eT�X{Z\�����i��P��ـ��E�<��;��ϟ���E(u�X�(�n�q%�n*���WL��`f����{;�N��BiQ3%rjn��ݟyXm��/���� ͭ����d���#�%RG`_����{L�fd���w=��נ1{�uU5"��㓽Oչ�`fֵd�ߧuXo^`��ɤM@��**��M�� ��N�`oe�f%�;y8�S��S�C���]}޹W_}��Y}����MFF#2��oe�`u�y�u=s`{k����^��dd������rWf��l�JgK::v�]<�2�r��cSlj�?�;���T�BJj��UK�{�~���́�>�`{��;�y��G�P#���'zZKc��M�UȈH�-��R���V[ם��kyI�T��UI*[#^٘���z)%�7����\�
&d�Md��7��_Rm�.��6����\l=�c2HD⑩\�#�=��v�����6gJ=�@Z�I3.����   ����   Xi"� t$` q�  �A:�.ٍ�� ��m� � � �b۶�ĽN�����ʗ{f�WcLǖ����u���&�e��,�W(�b��j� k�8[F�eGl��[VЪ dLq<������)F2>9X[��U�m�lc���f���ǽ���w��9��$䟔�H�A��y����y��yV����u���N�
nl�z"��J���ܥ�������n)Ȫ��Q��WR��<��U�b�I���g��,N�<� �a�iP"&��u%Y���,����*�IQ�ɥ���������#�H�u$�zN�1qs*����ߋ����>O\�wkKx1�%B���R��F�7{�7��j���0�=��3=�|�8�R�� �u��J�������i`>�~ym������U@V-�\�;YK*��NkX�[�4��3�Vͪ�b\9ڭ��K�"&f,��R�z�8P����y�eX�3D5�t�UD�v΂��ɧ0P��2�$F��C���{�����Ն?eL,�3�B'�J�T��}�� �=s�=Ļ��`ov�r����UMH�(�RS�އ�%��o�;��`w�֝�l/;����d�&�b�"�9%X[��xX	%�d���f�zk~y6��sa%7$����HI)�k��he�e&���<sM�i�+f[6"SD�ij�')O..*Uـw�L�u��>]nl-��/͕���}㢆�R7*T,�� �>wE�����d�B�V��\��*�T���>]nl��za�(.�B"!�(���@�=Bްl#���а�#4�hch/uvMR�9;'DƵ�m-��aa��F��2���2�(�� ��_�� Z 'iw֛0��� {)QAw��A�f�c^oon0bF�akI;��u���b1$�H�ر�a]�JH�#�<P����t�&f���h`%���JK)2y���+:�zݖ��h��q�	��S��8"qQ=�S�UX�i�C�G��n�P:v8(lENk��z6�M,�I)92Aޙ�ou��w�%)R"ff�l<���`w�L�A��y�PWoḿ��
���R��,͓�����<���gJ�~|��ʡgH\�-���t Svu�����[�.�ä%]c�k���upԮUHX���H��Vl��d�$����}���USR!
8Ԕ�w�|����v��>����C�o0M�ɤD��J�y����@{�:Q�c�;����F�P�wt�r�ԪJ�{3g��s��@c��PE/���Zf� ����������`b��]��Cn)�*����w�q3'|���@{�:P3$�~����l%�l�[:i� 9p5N~'{{t����^]rV��t�5�}����/��BMuV����s`}��V}�kOr"1@y｝��l��&�ܦU7�����߫���D�:V;��qn|�����T̕��X{�ʋ@��� �r�3j��W���3�B'�J�T��ۛ�b
^��ތנ�#ϕ��<�USR!
m]+�r}��v��7�D���N�no]�L҆ffL�1���   �p���   m�MV�n�i. $�h� @�A� �9���` mm�b�]�UUb�G3G�;;��$q|�QeD#�R���i
�bڶ�����V`�]+*IREY��i�!^&��*/I�ڱ�˚"d��.��6	���4h��Q�nwu.1%'ee;��]��)@[��E��i]*�����YT�,����\��YrE!Q��TE#�U��ɱ�}�bmkϹs�ޠ����P�I@k�9U5ˉ���u �r��^`.�6r����z��XqHܩP�>�����tP��� ��t�=�__�]�H!v�;����נ=�2ܔ��,�������g\�(�yqDL�M�#g����i`=z����K��~�����U:B��[+D�`R�n�8�mp�X�ݷK��Aj��$��ۣ�LyA���ݦX^���մ���r3����v�3Y�B'�J�T���f���Q�B�F��Gk�_����mX��v�za`y{�jD!G����y�(��z��2�Nɘ��٥������ ��#u�TE#�U�ݞ�>���X�Z��Q��s`?�%���T�.&��Xu%ݦX^����v�>~ɖ���UY�S�J��@Al)e,��9L�9����izv�#a�\�ڮ���|wbAj���%QT�MM��ـ|�����>us�>�L-����#�(�N�O���m\��]�=�1٭�d���z�>H�	�(|&&R�D��}u�K�;�r���~ܰQ�Xe&	 � �"�"	���H��"f(�&������a�������H�bb#�a%����><2gI>l>v�cϽ�@{��je"����}{�4�"�z���nl?r"�֬�CC���TU(���Qa�kט˭ͥ�Kg������=�l�}}�@�$R��R���M�2�6�hVd�����@JЫ�I�6�b�(�RUT�@��v���e{�z��̻��h+77� �źH�D1UH�T����""���v�`y�^`.�7���m�o
�R�-T.��{&��z� �u��;��V�;��IUIT��`=z� �u��;��V%��@5p��'j�=Ϸ�ʺ��=^�.LPA*jk0�[����V�za`nnoz�Y�Jc�HDIU"6�+E���,I�Z�ż��LWP��I\��m��)U7����{*�7�I��5�y��L�ٶ��T�a�}�&d�T|�� ��L�z� �u��5ovl�s\ٙ%<��B�h�������;����V�~��4�5f��TԈB��UL�b�\{��{[�M�!6����֖���y��-!�=�)�����UTP
�sb�N�z2t�;�z�>wE���wO��k�   	 -��@   -hM$kp�� d(  ���@6m�� )m�m ���q���l�� z��w��٘��3^H��4r��g�a�ꫬkM��3�E�H0*�d-Ĵ@m�G9�˹X�hh�H�9wB��b��rr���6��'�g}'_c��j:�Iu������}���7'+�{骛`�@ֲ�M:�Re����$�i����خp��mh��#��w�s�7�_�"#��y�|����� ջu`g����Cn)�*����67�ڰ<�U�}?L-�{�<{��J2�17`y�(}͊�=������%����L�T%35S��9!4ۛԍڦXo^`5��s`w��je"�)Ⱥ��{�4��j���C^V�Ձ�=�`|���IURE JP���SZV�f��v�}�n�&�:b&�f1u�;[I$�N*�R�U!�7w7���.|�5��ٱL�X���Ҁ՚��!��!IMI*�z�۵v���p�����f��v��z� 4�l�JjD��IV<�U����,����{�67��a��cl&��*r�+���~�y��X�y�������.�9���W�$�U)T��`6��q��o�?��ڰ>���./c��P�I��"�J�mR��bGH�M�į	Cj&�K��Դ��Dq�#�(�N�K�?nՃyY��ZX�y�`���M	D�D�P��N�N�{�����tz�; �8D�*b�Q�np�v�t��޻>mv�bHK�|t���	�|��g�nw���<��b�=�5͙�SʙQSɚ��m���.�6(K�eZ&&���wl1}�uU5 ���UN�.�6vWvl�ݽ02n�`�����U��vm5�@&\�z:DC;i۵k��u,rdu�^�[�,�T�%1����H��VXǯ0�[����6�7�r(떩]��@��i}\�L����>]nf�j����@n�ƫ�S(	9R�`n�os�y�V]�X��VfL,1��8���@�R�z�r!vwޛ�ܖ���kXy�r;��F�5�2A�
�i\aq��(]�7�iYCi���$_{7�4+8֠�j�T��5n���{Z���ޯ{0�[������l8�J�l�Ƞ�n�F�E�`�i]3H
lB�e�mњ���⺜�D#�K��j�6� �u��p[�V��0̒8�jW*H��kkw{ߙ&fR��&My��9�:(z3^�32lZ����TԔ��j]ܗށ矿U��wf����ŉN��8�U%5"d��UU6�G������֬�wف�DE�v�ޛ~�J���Lĩ����\��7f��ْ��r'��߯�ޚ����U�����?������h���]_���W��g��*���H�e�q���ֱT]����<�DL�Eu"�b�
H*�0"��J��"���0`UFBa����bH
A,@ I(*�
�,��+B*�B � !n�{�5  ��(�̪ P((A
 ��"�C$��U"PPH�L�PЩ
P P���R��P4�
2! (2� �
�� rG�_����ivN��޿������(�4
����n�?����y���1z?~(@ � ᯿�p_�ve
/���̜_���㤫�����w�W����=�N���#�?�[���οo�������x ���w��A?���AEEW}�**�ˇ�S�����a����؟�?h|����������Q����?���i��EW��ǰ����_5o���×�?���p��z���5���������s=f*"������~�=��k�gZU��=kI�Rd��"! I(	0�"2	
0�#H#B�������*�"�" �� D �"( � �R""�
$H@�	@)
R�D��*$@)$��2�H
B@)���
B
J�) @)) ����� ������HJ)	���
$�A*$ʉ$����K ����!������2�,)	!,�	HD� K!BA$$�� �� ,�"�! �$ #!($�!	A)$� @HA H@H����$	�(�0�J� Hʤ	"��)"@�
,�$$(�$ �$��$��!
!@($�� @�!+!(H�!"B�BL��ي�J��) �$H�"HB$�(�$�@�!(J��#"@0�) $!(B2$@��� �$# B�$�J� �$J J(@�
H������ � ��*)*�J*��J�����0�
2������(���,+,!,	"@��
�0�� @�*��!0,�(H�, 0�`p�e�dR�IFP$YT� FU�IV@HU Y��aD�FE`XQ�eV�%Q��` Y%��@P� Y�bfE_ @qDHQ!@�D	�eeaV$P�	RPY�($UZ"&`B�XT�!�IX�%VdH�%	Y��E"UR`F%T�F`RD%�G^g"_��O���������P_աDCN���������?�~��z��i��vtj?o������Y��'�_��MG��"���a������4 �����?�xY��r�O��Q����D�4���i������a�����������_�**��\�@ ��o��9�?������~���l�
��?�����ӌ�4��vw�o��EEW���f�?�,7��aqQU��G��y�_��O?��^�o�8���1���?������G[4��l��������G�������5|#����������� ����?���k�t (ݬO>?���y��{���?��?��?D�3������g?���y�oG��EV����������AQU��^�� ���W�����^����= ��o���Ϧ�����~��o�R�_���_����Ė��b�VO������� ����{�����pI����?Y�����F��?���PF�W'���������?����/�z�����B��������3���� Q�|>�QQU���?o�D6k��_�|����o?�������x���o�����
�2��W���^�����9�>���    h �   � P    @�  B� < �
�    T����UJH�D�$��"�
R�*RB���Q ��UE
�� PD���K   $(J �c ����f�����=n3V�� ���y�k��Wj�s�;�� �>�|���S�׀ //&����M����Mr|��}�w�nmҷ���W� �Rݟ/�����6_Y� ��Q@ �R��M� � �  � &��À  P@ &� 
 �� � �   �@)� �Q��� (��: P    �  �cJ J �  3   �@PH�� `Ae�u+�.c������3�^�#�}���׶�k�nM^�w�R�� ���yn����x �o}����jWw� �ҧ,T����g]�OiV� ޼k����o痹�wI�����  U (	Mdl�Ys�{����^��s����ڷ���P���O'���y5��]zyw�Wǀr�-�M�w_ ���+˓N��>�y�K���=�϶��=i�ӭ���)g{�}��7��y=v�oW��||�T@( (� >�W�Y�۾���wo���9:����gzӓ�m����Ϲ�����z]� ���t�Ů� t��v��K�� Δ��Z��Y�=�s���m/m��N;���mqd���|'}�_c�    ����)R�h0�S�H�7�R� F��=U*S�z�  =��#�TH  *�J=�R�   �jJJ��O�;���?���?��N�jO��>��}��Ш"��]���A]����!PEW����*��*��TU8�w��?{���\��̼�Ø���ٜ)�4�.�0��cL5�Cfr�0#\���3��I
a�CF)č0�6C`��5���L��y�q4q��� �I{��]���j�����Գ�xxx§Ν�� ��H�����$"�h�<�M`�S7���!)�55�8hv����m�xn0��8��0&��4�ǁ1LA0ѣp�9�7��.��@���j6%c �a V��`P	#"��Hb�CH��3f�J]y��rx}8�&�_�Cl���i�S�o�0m�	�>h���5��хM$��8��5�y�e�1	]o�������.�j`˗4]윓�f��]k���.����%�3D���y�<᥅�CF��y���IE׿!�9�!f/@�W�f_�o~y��I�x� B�7P�ip�$�6ō0!�$�k�"��� ��8���܌qp��ى�.x����I#� �c�$H�pa�gĹ���BF�X�@)A��@J� ���i�5�g6eߙ���n�/�����! �:G���kҎ���>_��HS� \������[���a\5����	
d)����HY��ׄh����i����B����8���u�xl�X�ɦ������>o�{��9��q���kT�{~ߞ�}7
�ё�@1cB�+D#�4�O�C��DV3�����1�.ߓ��ы�K�]�����MӁ��VoÞF�a��Ì�:J0��@��F����ńs��}����f�?�R4p�F�ȁ>��Xc_ ����ɷ�K�y��%=H�!e��=<1ӷ@��_R˭���6O!�r�P�F�JM����79tB[tR�p#p�ˆ�1�ʍv���F�h�
���F8f|( s��8�A�b� ��a��_��7�5�/�y淣

W4�$��T���M1��J�
������i	}�d�K�|��s��w)K��|H���=Hl�5�&~Nf�̸>���:`��"~p�-��dB����{}׺3$!�.�C���ÁaR�h�m��s!��`R��l�
f��Å8�ƘM;!��i�a4l�(��n.1.ac��JS0͙��a�v�q�p4�6c�X�5�ه
��p�v��1ц��3D	!0֮���7�/���LJ�@bD�ư֡ra�y0�Ɔ4�!��9�.�f�f��dt1���7�24�&��Nl��L�S{�p�3w�<�9�p�0c\3	��Y#J�f�É��l]FzzL5�S|���f��������|s�4����/��		5i�9	���4h�/ �Xe��o�,��4l���4$�#L5�M|��B淹xNsP��F��k�2�0<3|�!��O��ܚ�;asz�9�{�a��a��	牤��4�H�Ą��i`L�8b����i�.�>=��7����k�r�E�,�>0�V�2!�I����4ɛ8O|�aK���r� �a���<�ֽֈ[��[�Dl�Q���[�^�$J�ȯ([�*�o�R�R���&�ڝ�\�����l��{��F�M�C�D"B�*"9�kf�V��F�O��jP��p��捛8Jp���Wf�HpesA��B�����h۳�hF��kgc�bƀ�F��"�#
᳆�O�F��߾x;4�NĖL4=W;xH,��gX0�4l��qѰ��3[�l4l6�H��[8;"�[�F40Ѿ	.:M��h���$!8P�g�.�y�-D)T�dD
�-�v�)��T�ĸB�6m�cp��F�7�D���/����ѾJ��-�HH5"I���T�q�M�<�x�VD�,l�Ě��8��.��B��[�^d#
f]a�8��h!��$.0������fMa��)�t��<I	La��0����F�p$D�ч��,�!��#�ґ��@���,�0�h��
�t�|�H0%a���W�,�]3g'!���1�w��14�&k.�o��M,+��¼�l�8�ư�4g)Œ\.����Ҙi��8b���<9���Ȓ-�@���HIH�2%"H��ė��3$��RHH�̅��#H�\�e�S	#d�����ӛt � ��E�>Ҟ�۲��A��1h�h@i �d���a�6�R����SY��y�4s���B@k&���|������,ddZ���y�4뜄�֬�������5�P�vE�����~�79~���:
0 �S��
�:���2��B7M�Ԕ�dZ�.��Z�0�j4调S!`��3c2M5ZBɅ�#H�D��o_{�:��DnE��D�s[������0��*�EHX�PH��d(�D�[�6�S�Jh����B��B�j�i� �D}b!P�AX��ٯ5,�z|��S�/=��O�׳̾ۻtsÒ��� 0�.�o���D ��[�Ņ�[<5���H�5�gx$
��g��sZw�;<OY3Ro��׆�T#ILֶk�|BY3FӁ�׉$)���pߞ�)$�i���f�FT�hپ�
B�a���t�	JX�в=�6U���*�n�us�_��_��TZ�_�W�Bj"[���a���+��7
�g���m���(秙�Mzxy�"��׾��5,��сXf��-��㠃Sj�!VS5�=B\&����I
B�:V�8�t�G$$ae��3�@�i���vJp"�G��������<���~������vows�w�B�Z����-T��"!�z�+���x_i��5�[)�h< ��Ȣ���מ��C�I�!％�k�pc='#S$�A
a�1�6��tm%ÞK�y�==}��#㆖I �4E#"Մ�u�@�h6a���3p�Fc��%0���G��]&����fÐ�n7tn�`rA���8a���%1�x[#�P�na7�)��.��9�p`�4a�ُ�S�c
�4�o��Ѵ�o5���֙��/��&�hۜ�<4oa�d,h0�"V���槳ئIZ_sg�>�|8p�E#��p��t�h��P�Hx`��.y��c0ӆ�9&�h�Jq%0�[�zx���d��^2�jk|$�6h��B��6Hp�<�!sF�5��4����&�<%�!K���a��#sRy��T��Ǆ���uꐸ{>D��A�e��7�>�̻%���":�	������a}cT�B%B1$����d���{���Յ�D ���ݞF��s�4)��z��4L�xJ�BHBM$jE��Ad�c$�	2@	�XD$5�$L��jC��<}=6F��Jx���6q�:&��jz�jX��bJFJXF8�rc�`�3��D�@�������p���z�^���Vz���{�Cŉ����F�8h�{����J�	�p�D�iٳ��%�7�܃	
L���f�4�Mvm8���"��8g�珡�	�X��b�dߊ�
�R�^�3!�kȁ8�B���f�9�"�"��L�
f��LѾ��8{	cY ռ�@�XU"A"Ő�Y�3�rk�)��MGk*MjSy�XɢL�Ԝ ��"lXV`�X�&�H%$!��lbT�h��������І&���5#���� a� ����a���Ѷqa �!���C"h�3R3o��I�ǀ@�
C1����0��8	�4�g-p&���Ǆp�M�)�%q��9805
3	&�3|*I���8^�M�p|d�0&�s�4$�r�M��B�	���
5�wʛH�.��a!�h��(�s�}5�k@            $                                       ���   ڏ��3K�隝�*[����0��-RY���
�	VVV���e�g�N椞Ƹ�sV��$�W[R$�aV� H:	�  *�����l.�WR� 0i
3E����*v�\u�@�����B!SM�m6�"�mH*]��r�6�XUj�6�:D�:��;&����WPsJ���lm�              m�0               �       �      �`                                                               m��  �                                                                      ��m��                 8       @               �&	�6ʶ1k�i�j�����:�z�e��%��l�vk��j��}� �Y���R���h��m���Tp�vv.�@O��t��Z��U2H��J����\���S^��ݙ��n��)�[���� l8�_&�I���j���rt���q�$���ݾ��#�'սM��5h�Uʶ�
UN�.�\u�N�� �� [A'6n�nʹ�"մH �(�V�mu�1t T��ݳ����\]#@ h�H�Rn�i8�r�`��Pj��n\��g�������Ei�� �[�� Im��u[x 6��p��u��ڠ��^YP[V��l�٤��m�Am��*յp��+J�M�uI�C�Ŵ�3GP�g���rL�T�����E�`�$n����H �C4�l�N��}����u�j�Kn� E���� ��@#�v�Eҩ����!-��� i�Y9pm�;r��l-*�*�T<vݦ���'m�Y� $n:]c���M�#D�Z��b 9tj�A�X�mH ̙6ؽh	���v��`j�Z4��-W��� 
kٰ+i$M�d��m%� Gm"�ex6.�h�[t�gk<�XΦڕj�M��^�6;�:�%�ɳ�	-����r@	��  u�HZm"�Ӷ�A��5-���]f�z�V�"�qm ����m��  �`$ �I�B�bn�4�l���+�(�9�v
�V��)Z���&��U8Cf#M*�N�L��J�=I.� X�r^���mv�K3 �i��������[�{�QZ��݋�������ɼvU�x���T4I{m� v�Y��E�˝�*�|��]�%V���i����݇�~���t���5�	���|��[�ʩ-���/t�T�c�P�j���a�{Q�0R��[�O�tk���R*D6�m�ϭ�~-�n��o@P���qu
�Ѹ���zΧmQ���&��m� p�"Nε�l�-�lݴ�Ѷ�  	��I�ϫ[d���aΞ���J�!����J�\H�l!��VV����j�r���l��D��I���m���f����h��^��ۡi�ftt��9¬uUP%�Q��֓WUl�k<���c�VV�\=����m�`�؎t<2ݷX.��wk6qA�ԫ!�@Rqv�F�����c��8�u�@������;N��ntt�	����[�9��:g6��U���BiI����ʵt�^Z�����ГT�@ʚ�vI��/R�mJ�T��l�0ʯ:i�m��	tY.��Ź��t���m��-�I�z�	���XI��b�Ԑ�cjy%C�Z���5pq!;�dE��Q�6%m����3�:�ۛɮܓ�C�ku����ۉ6_P  G!���WiUv`k��^iI�j���°h�j��⣛Er��]�ϙ��?�.�=��gj�]��)�/6ۈ���ҭT��-�ݭʶL�g-���m�V�C��傐Ux'�dfWoM��[iSn&+fYd�.��i�f�  3�2�	 q�@.���yɤ%Zϖ��QS� 2 �� ���-�mm��}e�U�"Sm���       g��+/UR�(s.6�����ul
p;*�Qƫ�[��&�6�S�"�P�uĻs̰U+;m�zu���rA�����v\-�Y(�oR@�iv�B�Oj�<�1Α:ͷA�+�r�@UJ��\�ی(b����卸�`%^���c`ح�fҼʁnR���O@S�8Un֕櫥�`*��Y�Uj�ڸz�ŵ5ͤp}o�|mm�S0R����H� {"]�t��5�/+�3�
t��8�]��ڵ�[��.�:5mhɭn�,Y�cI��t�vZ-�"E��Ƚ��I	�eƍ�D/z�
��J3fJ$M��V����P �Ĳ���m�$f�
�����]�Y����UK�KJ�;O*��M��6�ip�Kne��m�I'm'sj��]�y�,1��l9�a�p��l����fͰ��b�&�g�(�n��	V��+� ���bA�m�"d`*�.� 86+�uUJ[-cɶ2���mA�Ҭ��U������+m�m ��	�� p���r����m�p�ے�HחY�����lMeߏ�|$'@6��ܶ�H�dt�m^�����ޢ��S �kҦiP*�C��9�M�'s�N�#
�U�8{]2�����[@-��&��`v�m6�-6$�i�7'���f�Vm�*�.� l�KJ�y\��!5m:�ݪ�EHI�字��(�X*U�@	�6���c������Q��N-ֹ�vZ��6��U���`-6	q؁�-�[�n�	U��i�K(	 �kh  �`�      4.�Vձ�8��L�  sӤKYj�L�92HE��PA�!�����t�4����:吽�� ��t��$�7knN�  n2'C˳;�^��ڨ   �m�  m�D� H[�� i1���ڦ�
]Ζ�W����j�Vy��ޚ��Mt���0T� k� �    @ 	,���Fl٭�8�ֽ�8�ֲ��wn��F��� Hu�i%(lWA� �U]T�V�kZ@ٔݵӱ�`])m��c �]瞢RݕڰVҬ�@5MK	!�*�t q�U ��am| h  6���v�AmCz޹V�&
ZR[�|7�>smUU*���p��,��UBY�R�)��l֦k@p��9���o�k�n9l��  �lņ���'�N�i����pk4�BA�nͻ U��!��I[ڙ�ͫb�I�r�l ��'ku��l6l�q�R�P*���;�kj� .��anrLT��k�/m�V���v��m�$�j�[v� ڨ Ը��v{e|�UE��[-�6�6  ���M�      t�'���i��[t��2����*�mPUR@         ��N��H�q���(8��		�m����ii$�c���>wϕU�J�Ӷ$�` 1��mQɜ(T*�[5UUP\i��_@�]�e�m�P�5�̪�ҺFy��,���.n@�C�O+WJD���7mPY�N"�:$ڵ��m� +Z�P�U���U!��;���� [smm�\��l �;��m� ����`�6�����k�ؠ)]�R&�%�)j���8ؕU�W�ZU�ڵM/r�U�J�@U\V�ݐ�j^����)���Ij�	��]/T젌��"@mK���,��mJ�T���%Z�U���U��`:]L�A�J�����St���ut�*��um|��#���(v�A]���Bz^�c��J�2��G	�*�mF���Z����L�0�[j��e�u	�؄�:@;ol��h�5sԬpU/l�UU"���`�e6�f8�i.-J��vQ�s�GY�TnR����2tUr&{*mu�*�]t��W=�5`s��		c�V5��VڤP�-���Z۸�s�,��Q�3��햶�r�uN�I�oTk6�nZ��]�烶D]=��RɺѴ��j�1�wnW�
��`*���Vv:
�(�bt�g���v^ګ������6��&�$���I$e{e��M���]!������BF��7m�:H�$ڦ�-��k��GkW��I m��L6Ͳ�U�@��VV�l�][[m�UѰ�0�m2m�$���$|[rUR� �7 �[U�U��6�^m��q��8U6mГY�M]jL������*��  ���҂�D?�P��*��@@��?ҩTw�G�QB�� A�M��(�8��"�Q �M*�B����	!!	���#$b@�'�'�&�>8 1�Ҳ)O�x!G�T�#�p���/��	#$F�!a- �HIY�B�D�!'���=E� h� �	 � :U\D( �"|�b@"(�⢘*��A���ʿh��*����GB��A���O����l��"@*��P�W�C& �
����4gE�H%�!$$�� ��`���$d!�1_ �"|�I$Z��~b�� !HE� 1b0��a$�D�=TV�Ń�'�� (�' �E>�-�Bz�$"��>��B	��h���S�� :�@Z�!�PQ�>(0P*��E��b�D�TL
��!����������"�� �*1Q�
�^���?S�  ��       �a�g4ގjq3BW�u����LŲ�KC����f\��6�   m� $             ඀             /�  #�   ��ۣZ�d��F��D���QC[w:s�0Љ�Itҏ��\�Gf��N��uC���7<�� ��lX����v��-���=�f&�����-����G:U��v�puq�赊� ���m;�'kks�8�en��u�ٝ$��u�m�I� N�ni,�M$�դpԶl;
R�5�9�����.n�z�����tbz#��������Uj^��t�_JH�q;�n7GW<��T�ZL��ZH't���t�I�]���� �q�Pٻ8e[lGh�6*�õ���g��m�2nΧ��y�[��UV+����a�7m���PsM��x�����tv}2��<�݃�5C�jS�tÀ�e�:M��v�j���F��g�3����v�J[�Z���m�ڞ���uSx�R`w9���iv35�{Y��)��7l�1ל�*^�ͪy@y6��x�t�ۗV�V�m��a�9�6�v�D!l�-���]n������˻9	�^1�Y.��^ۖJ]��E�` ʼ4��q�["��g�ul誮ں^R��j��&� ���]�����gv��lp��!6���۰$!���/ f-T�����:�팠�n�t�:�����ݑ^�-�r�!��v9���N��s*�mT�z�KPSre.���ZQΊꞷ��魃��6�\r�ric*ݲ���$���g�5�6�c��$rj�2s�܅ �� ��ٝ5���-W��,w�����M烴pC.��p�s�m�D��g`K0Ĕ�p��+��z�!�X�ѣ��<!=s��8�z�'�!�m���,���.�5�{E ��^��*�­��=@&��!�
#A��� t#�k-�kZֵ�e�Mq���ˁ�@   �[/e�tt��5�ׇE�s�vR�3ڶ�7�kBpr��.ܷc`^����+eG���I��k�v�Ů[$�����t��8�ڔ��GQ�爐ˎ��3��s۶�iS��Ή��֗�F`�MRn�X* ����a�[d	WFe�F��m�6���D,E�"�b1�ْ���qw��:�ʫ����� 㲛��7#����n����g�bX���o,�8d/���;ޙ �}���}V��-K��"i7y�v�`Yk���`Y���ژ�yδLp$S$m���{���$������W�$��v�J�L�Z�!Bx�s<�$�;cԒW�j�Ē]n�RI^��y�I,FwS&6F�F�F�z�J�-^x�K��jI+�|�<I%���$�ν�m�l���D ��C�QW]����Nm=��L'�VbS:7]�l��JH8�&Bqy�I+n�RI^��y�I*�RI_e��I{�UvL��2b�$ԐԒW���x�~���~�$��=I%}��<I%m�jI/3��ߒ4��%�E&y�I*�RI_e����f~�͵��l5$����y�I^b�I�Rd�̎H�$��Z��$��a�$�u�<�$_�g���C�z������%m|4�VK�}�I+����W�j�䑻��]����N�ڀ83��2�Hkp6�{N����%�ꃉ4�yd�6�] �nCRI^��y�I*�RI_e��Iu�I%_�s�L���!�&�y�I)����W�j��R��I%d�g�$��e�d��ۀ�H܏RI_e������oSv�~,��߸s��}Ͼ�� ����;��ζ�L1����}�5$����y�I.vǩ$����$��*�&Hԙ1d�ԒW���x�Jm��$��Z��$����I{,�~�7�,����t�eH�t��(K���z��v��q{:���ՙ�$W~~ ��{ZI+�}�I)kᤒ�_��K���2I�Rd�̎H�$��Z��$����IY/���$����I}��~��cI�����Ē]n�RI^��y�������U��z�K�|��$��u�c�"�26��ԒW���x�K���I+����[TOQ"� �@����jI*�3�jdD�q�73�IM������W�$���I+%�>� ��}��l��hց�̯�z6�i�q��,W\vM@�ĺ�/M��΍���n��F�a#r=I%}��<I%��5$��g�$��lz�K�͢i��8Ʉ�$��ĒR��I%d�g�$��뽭$��Z��$��eU��"�&,�C��J�_3�Izu�֒J��_|�JZ�i$��d���2vH��� ?���? �����$����J�~ϾI)7���w$-h�rY��n�o�k�9m�TC>�y��m�����-����f��P~��o5�ۓfmՖ���p    �][5�Mԣqlu�P�f�@���O�Ǵv>wB��qϞz/�N���V����P
�&{3���cNJ7����q��F��l�ܺ��3��r��LqO���j9{p�f�5�t�Y�ڳ��Ev8�����E��:��t晵�\�=�ܓ�ji��m���rD�F�k����$�{��3��V�]���7c���n��2t*+�����rnm�A��խe�����I�1�� }���f�J�~ϾI%��{ZI+�}�IMܛZ&7�1��NCRI^��y�����?6�����$��>�y�I.�a�$���u���6$��<I%�]qjI+�y�I.�a�$�u�<�$��gS,����8�ԒW�j�Ē]n�RI^��y�I/z�RI^��;"�qǂ[��IK_$����|�Kҽ��I__~�����}��UY�7n�PeA�s��.���Z\�c��O<F�nqf�����1d�ԒW���x�K޺�ԒW�j��ZI_��jI/s����'I�2��G9m��~�j�x��P
Р���
H�4C 4Il����R��I%d�g�$���U��@�ɉ�IZ�J�-^x�K��jI+�|�<I%�]qjI/j_�'148�$#��Iu�I%{���$��-I%}��<I.o9։��QLj&��������Ü�ު�{�y�����{��r��[�ԒW=��8FH���d�@�P�Z�jSN��^z����8��ق�ogW��]�$ȉ�8�ě��$��\z�J�v�x�K��jI+�|�<I*��ǋ$i�l#�8�$���<�$�[�ԒW���x�Kޕǩ$�gj��qǂoS�����oSv�~�߸s���DUt������$����y�I/pʫْE&LY��ᤒ�_��Izu�֒J��}�I.�a�$��rѷ�N4�cQI�x�Kҽ��I_WO�I%-|4�VK�}��_}]�~ʶ���\<O�Wl�9<7���2�ۥTݹK�}�;R��1]q����$��t��R��I%d�g���}�~�� �;��=��p�/5�ߟ$���I+%�>�$��WkI%}]<�$���Z&7E0pi9I%{����$��ZI+����$����J��Z�1�1���x���f7n��ԭ�����-�����ݷH� �H �3?O��^���x�U�2�,����$���I_WO�I%-|4�VK�}�I)/�� ?����_���Xn8Ԓwchu�S��;�ϩ��V�<���Ӯ�ś�q�����$��v�J�_3�IwJ�ԒW۴�Ē^�W�$�L��	HjI+�|�<�?6Ҷ|�Ԓ_w���$��I%�{���"q��梓>�$����I+����$����J�~�������u�uù�G�?{��k��q���̾�&fe���tDB�}�^�>�/�bs��X���u�4�w4���/�S@��e�Ҹ�I�z�Z:ꦑ���H��  v�  �S��R�iղ@ �r��������%�z�<;.;#<����ǰ\p�R)��ޥ��l�z�fk�p��x������ъ���y�;]���s�;*Q��n�fk;!���(Pg\����v�$2�-�ew9^��
��D/[rpR)t�{V�:p�\,�k.[p֌�"� v8Moz��u����]y.�����׸,���c��]vԼ��q����5�lEٳ���o����x�%����0	e�G�M��Z�7WE���� kl���Q2v���^ �^,exM�)Wu5aJ��|s�����^0	m9�ftCv#� ��4>J�~�����m&�}���ʻ2H�Ɋ���`Y+�-�0/�Q�K/=��������J��ݪ�:����[�=��]v{��%#��T�nDw.K���+C �_�r��-�0/�Q�K/0,��xk���ɉ�bf8�4�������DF#��EW�y�d���������Ÿ����7�`��%x�%�����*��Z&7E0yNM�]�V�Xר�%��Y6��옣�������z��h^�@��s@�T��'�ؒ��L����g���\Y���vq�=�[q�u�<��6��ݛӮ�W;,����$��/�S@:��+h���u�$������k�x�x���X�gD(�#*��2H�ɑ�I�&���nh�����~O7�C�Ny� @'9� �їg�^���!f����aq-�K0�-K/���Cd��<�9�¨#tS�H!���v�apsU�"bi�:BR�aR���Z�)��
�L�M@��m�Y`�T�R��kR�"I��s�$H���9��84�E�g�J��F1+u�bLRS	"�[�XX�L��!*º�J2@d�Q���D�r�h!YIFRT��%m�a�f���Q#�Ť�!
B��e��8��&Ң�P��U<E���\P<<X�� ��J��T@��͠���{7$���@�=�F�AƓ�_��L�9[F���F,���W�So���[��Zi�ư/�Q�K/0,��+h�1r+U�6�?ͨ��x��÷>�7^�06�5u'bv竷u˷/Z�A�C�˛�� �4�Y�^빠r������w��@�\�才�QLF��@�W����/�Q�K/?�ď�E����G1���_}�����f�{���=2�`�F�����?;f k�x�x�)5
�!" ��A�� �CH�89��c��@��$I#�0p�	e��ex���kzvp{� �iVլ7j7�OF�i�v���F��v�F,F[�v��sq���I]t���7���6[e`����H�^�v}���8�p��QI�+h���0	e���`Xj�n���97Wo���F,���W����"Կ\NccpY�4�Y�^빠r��@��M��u�2L"�WS5w�=׋ ���w�޾0�{��krO4����T��EV)A�D�_���4 ݤ�ər*n��� �l  :����a9VH��t��N9:�WO�-����-��]�Vq1u#և��-�&/L��٭m�n�;h7IZwqɺݺ�0H�,U/*���F�A�<FL���%ݽ�?.���&ɝ��a�R6�Z;��6v!E������kv���j��,��n��=�MM���'EaRK�uWdݖ)AWg�D$�D$�?%p�J�k��n3���*�ys�1���7��[�ny�V�*�֫,�V��d�/ 绊��� 5��X��c�4�<��z��h^�@��s@�m�{WcD�8�Swx`��%x���k�����$mI�#��RM�]���z��h^�@�=�F�AƓ�_�nn���+ �B]��~ |���w4��+Z�ly�� q��s�b������ۆ�ۘ3�����%��o/<HD,mG�_l��u�4�w4V��"Կ\NccpY$NC@:��ߝ=#H�bB�B@�� �1b�$%JZ��(J�`��:��`{����3�?f$|�W�Dd�8�#Iɠ}oۚV�Xר�-��Y6���q��*��@��M ���/u��=�8�,s����A���`��%x���k �fSwK6��"S�wTAΑ*��N],S{:�j�v:��qi���jf{l��`%��J�����0"��Y#jL���5$�/u�߿~�ٙ�wqXo_�]���eV]�u3V\�M���6[e`�م��&�B H��
"-%!f��?6�`J��J���3*�n��J)��� >��X
%�w�zN��5j���gp��`��I^0"����^���z����p��#��_����e�y�����;N���XZw]z�X��ɋ����nv���I^0"����^� ���=G�9֦H
H���r���~�l�kw�{u�΄�����9��X�I �o��@=�f��u��=]�z�al��8��Ln�n�=x�N�+T(��,�P�{/��*�b]d��2b�$��@���`����^� ���$EZ�`{2ɞ��s�k*:����#���m�O�[5���0]t�2���6����������W�So��x��F1�	�y�S@:����s@5�^tB��='t�r�����*웻0���=��a�BJd}�^���Wg:ЦI�����= �e���0:)��׀l�)�Tڻ$s�h��@󬦀[�h�x�Q�z��e������+]��MZ]t�		     9��ԑ�3�=����VٷL��)��[V6:ykp��Ϝ�|pR����ru�����Wp��W�D�0)�n:��n˶Ԕɣ*voY�1d��E�:��]��x��P4�CQd�n���s�&7Iڧa�#�,��i ܦ+c���}u����4c,sҮt]/ӛ�㞎z�w����>B�˩V�h�R���b+N��a7E;s�
�����.����<̊`�F��!$&��Y����^/�G������.���h��� �y�d�� ww�~�l߿$U�%~�6���HrM��s@l�?�B��IUo}�w׀~Z����Ɠ�_��L��?bW�&���|`z��'[�� l�u�T�Mݓ"������f������, m�h9�<x�����s&&ы%6:
WG2���[��me�]:H����2O��ۑ�s�x������~���s@:�O�x�����>W+��2L��F'&�<�߶l_� @Y ��V,��	U�T�x����I���MnI��?� ��o��#��+����9���X �����s�С$�P���� }�b�<�h��%]�Յ*V]�x�O��N >}x��X��}�^ڨ�}$�"�<�����f��g�}�x~��h�hV��7d�H8t77+�kl@�]s��Qs����vn�`+��4�>���楻$mI	����:��, m��m7=	/�s��<�|UUd��5e�\�լ m����$����Ӏ}�^�ot(S#eK���Jn�ue��p^��T)IBV�%�EN��X��/ �a��t��6\�]�(Je���5�b�m���~�]g�-�r���0cȞH'&��o�DBQ�IW�}�~�}��}f��{n��2D��%25 a!>h�E�wll[v�΃����o3؂�]��������t���d`�� >�{�ՠ���n��y�Ud�8BHM�M�t$�C�����`m��	)G݌�}$�"�<������M�o
d�|� �]Ӏo�L뻺����%]�%�������m7w%�"!��`�a�7����rO2��m�NA8E�)� ��M�ߺ�t� �}x��XS�uA4�F�u���t�i���_]�zt�v��J��sr<mR�FE��<RA#�4yڴ�w�{[�ߤ���Rq����.��s5w8 ޻Ι5�b����k�hvs�
d�7�'&��[��-�9�鶦l���<�m���
H�6	��z��=�j�z����}�� ����l�.�j+.�^�� �D(����� ��`z��A3lČH@'�O����K�p��(J1�
a�<B�'��$	,����0��ǁ�烤S^!�%�db��!���.�q$RZ�aB�A�	u�qhȑ��#H�|���#�!	&�KHR��Z��x;6£
���tD����%� �=a ��vx�	�T�%IB�B5`��eeBP��
(H�Z ��Psp :]Q�T�:9˚� !@��V�R5����|4֕!Z�!����� ɪ�ӈD�#�&�U�ﯞq�F�C�XR�IhJRZFx�w5��4��>h	s[�_F)uSF">�xB�&$(D ŉ
2����
¬����)
2��ӯ�:�_zuߏ��� 6� ����    ٭��6��AT�uv��h��������ص�y�Km��>}��m�      	             �m              )�   -�   
��i�9-�����c����aJxG;���m���X�5�y�u�L�M�t�&b�cOK�ʻ/kp��<v���ko��J�q�j���n�嬨S���@�J��#��.�L�ͅ흺g�n����)�u���嬠pt&�q���u���)���q��
���Pv�u�m��6f]��=� ��vq�4�X{$m��Ȥ��k�ۺ{Ng�e^��^ٕ��Dt!����|L�쉋�Zd�M���"�ڻ�6�tnշ	�QK�\�f���k��Rvt��\���]�M\����Qm)Lh���)a�0� �c��UV�������`Ѳ���:8v�ҳl�۰ �f��۳�-Eu��%n;Ƒ�8�sNCcX�m��Y�����9�g���⶞v�Inܦ��X���6�;`ojeA�.Ϝ�8N��m%�;`�qQ��R�i܎���UVq�&6�=����e盛u�H�X3���=[���^�i��vJd���D1�\0T�3Ek�m̀ �E��jW�흌�Q�୻i��S�6�YSn�G:�N��ɳuU@[*���wm����6��\���6>|�}���T�&I�io6���0[m'vζrl��9�kQ��S�K�lv�������n	��U��v�)���񐖠*�ܴ�v��&v���\�[u��gi��p/�����\n��u�7m�l�=o&6�H.xCp6����<�+lr�K�;$q������v����;��m�u�wn'��wO;����+�m�g��R�+���O&�3�?>6���;���M�y]���\�q�M�����.��Sv#Ռ�5�x��(��t�*��
���⨼<"�(  x +���O��kZ���]�����\�H  8  W4:svNŷ�p"��yy��c�O]��[����C��lb�����\ѭ�ݹ���XS��<��G<���}�[ڋh�nz"β�cy�;/6���]˦ں�D �g>L����nSN������*�+�챶$��c�%�v��r��xh���\�v��^��T��<&�YfjHc�K�53:� 9�I�yiV�a�<�I;��sI�Z�m��Ɛ�q�`�gH��3f��~�ܑ�Fn��e�_d��߻���bX�'�w�6��bX�%�~魧"X�%����nӑ,x��{��z��)V�x���{�7��bX�����r�bX�������bX�'�k��ND�,K��w[ND�,K������\֥�MWWZ�ND�,K��t�ӑ,K���w�iȖ�b^���iȖ%�b{�{�iȖ%�b}���:�]f�a�5��r%�`'�k��ND�,K��w[ND�,K߻�ND�,RĽ��5��Kı=2vv�3F����j�֮ӑ,KĽ���ӑ,K�~�xm9ı,K���[ND�,Kߵ�ݧ"X�%��;�u�e����n�F���2�Q����n{zttH�V�N�4�Q�v:w���}�d�z�.au3SV�Z�r%�bX�����r%�bX���Mm9ı,O~�{v��bX�%�~�bX�'�=��ܺ5�5���0�4m9ı,K���[NC09���1��cX��P�P��H���	ӆ��$�x�H��bw�{۴�Kı/{�u��Kı=����O� fDȖ'���~���kW5&jk4kiȖ%�b}�~�v��bX�%��w[ND�lK߻�ND�,K�ߺkiȖ%�bw�R}�j���a.��sWiȖ%�b_���iȖ%�b{�{�iȖ%�b_�ޚ�r%�b'�k��Noq�������}��J�g��W�w�Kı=����Kı/������bX�'�k��ND�,K�߻�����oq������~�*��v����tӷWq�Gv���;�x�����܈��.;_=�]S33w5�sSU�ֳFӑ,KĽ���m9ı,O~�ݻND�,K�ﻭ��@�y"X�'����ӑ,K��ٯ��Xf]f�a�˚�iȖ%�b{����r X�%�{���ӑ,K�����ӑ,K��o��9ı,OL�rW�5���[����Kı/~���r%�bX�}���r%�C�1F �}T@좤��ț����ND�,K�뿮ӑ,K�����Is���f�j涜�bY��"{�߼6��bX�'﻿��9ı,O~�ݻND�,���!s}p���!zM��m]��\ڪDլP�BO�˅���^��9��,K�}�m9ı,O>�xm97���{���v�����a���cs�UI�,����یq��{Nf��/Ok��kf����2�nӑ,K���}۴�Kı;���ӑ,K������9ı,N��yfӑ,K�捻���5�5��]2�WiȖ%�bw�ͧ ��bX�}���r%�bX����ͧ"X�%�����i� X�%��M[��Z̺��ۓZ�ӑ,K�����ӑ,K��w�m9�����>���9ı,O���m9ı,OO��2�&kD���j]kZ6��bY�D�D��yfӑ,K������Kı;���ӑ,K� P
*FDW�*U*�&}���r%�bX�}5�0���5�Z�iȖ%�b{����r%�bX~T������yı,O{���"X�%��~�,�r%�bX�����ܔ���#^�G� 0�ϳ���v
��WRu�ɒ��ێi�0۶Q=s�Oi�c��x�,K�ﻭ�"X�%�����"X�%��~�,�Ȗ%�b{���ڿ��$)!kO��k���eYd��AȖ%�by�{�i�(X�%��~�,�r%�bX����v��bX�%��w[NDı,K��>��ѭI��]d̙�6��bX�'}���iȖ%�by�۴�Kı/~���r%�bX��ߖB�B������M�%��XR�.f��r%�g�B �D����v��bX�%����ӑ,K��߻�iȖ%�!bw߻�6��bX�'�5'{�a�Ѭ�虗Z�ND�,K�ﻭ�"X�%�/���ND�,K���Y��Kı<�]��r%�bX�~��w����-�� %��hm��h �l  $�f�͜�d�#�<�T!����3�i:�:0��Ļ��;\���f1]֣i����n�)�8�#�kR9c��v�i�����`���nCl;qΎ���{���z����ú\�����U/ [u���^�i{�*�t-���F#v#I�Mog���ͥ�q��h�M�G�4�j�+j7��綗v�3�,�)�h�F� �q���8��ub	�Rn�|*�{��,K��p�r%�bX����ͧ"X�%����a��@Cșı/������bX�'�O߳/4f�K����֍�"X�%��~�,�rؖ%����iȖ%�b^��u��Kı<����r%�bX��k��aL�k4[�]jͧ"X�%����iȖ%�b_{�u��K�W"dO~��ND�,K�w�,�r%�bX���+�	�Vkf��j�9İľ���iȖ%�by����Kı>���ͧ"X�by����r%�bX��}��.sR[��f���kiȖ%�by����Kı>���ͧ"X�%����iȖ%�b_{�u��Kı)���L��ʶk��n3�n���p�끝oD�?>d��^y����:w_��|����V���ə�i�Kı;�rͧ"X�%��{�siȖ%�b_{�u�D�,K�~��"X�%��t}�[n����2L���iȖ%�by����r �G~�bdK�{�m9ı,O=��6��bX�'���Y��O���{��7�������=7L�.�Y���Kı/߻�[ND�,K�~��"X�E��L�߻��m9ı,Os��ͧ"X�%��O��ֵ�̺�.4��kiȖ%�by����Kı>���ͧ"X�%��{�siȖ%���3�����"X�%���������F��.��iȖ%�b}���ND�,K�C�}�ٴ�%�bX������"X�%��w�ӑ,K�����w㪪�vb3q�ۊ�h��׌;�����^c���\��v/Z#Ol-<r���s%�6��bX�'���ͧ"X�%�}���ӑ,K��߻�j"X�%���w�m9ı,O��醬՚�Y���fӑ,Kľ���i�~��L�b{�p�r%�bX����fӑ,K��=����Kı=����fsRL�u3SV浴�Kı<����r%�bX�{�yfӑ,t��. ���'����ND�,K�߻��"X�%�}=��ܺ5�5�����3Fӑ,K?
�P"w���ͧ"X�%��}�ٴ�Kı/����r%�`~EfD�����r%�bX�~��~���kW5&d�s5fӑ,K��=����Kı/����r%�bX�{�xm9ı,O����iȖ%�bS߾;33u*ѭb���Ť�%=��mM�t�S���69Ε�/4ϻ����O�/3��WL��ͧ"X�%�}���ӑ,K��߻�iȖ%�b}���ND�,K����ӑ,K�����Z�f[�3\ֵ��Kı<����r�"�2%�߻��m9ı,Os��ͧ"X�%�}���ӑ?1S�����j%�����̼њԗZ2���Z6��bX�'����ND�,K����ӑ,Kľ���iȖ%�by����Kı>�k��aK�k4[�]jͧ"X��`��=����ND�,K������Kı<����r%�`s�$�"�@JRAv��v��1 2'����ͧ"X�%���_�+�a��n��j�kY��Kı/����r%�bX�{�xm9ı,O����iȖ%�by����r%�bX������m:v�ӟ@��4:��ۀ�; ��n�SvIjL��]m��7�|̓9�Y.]S55nk[O"X�%�����iȖ%�b}���ND�,K�����?B)"dKĿ~��m9Ǎ�7���N��um,.[�{�7��bX�{�yfӐ� �DȖ'��fӑ,KĿ~��m9ı,O=��6���)��@ E5Q,N�h���K�j�̓.f��r%�bX�gfӑ,Kľ���iȖ%�by����Kı>���ͧ"X�%��MI�u�k4k5���.f�iȖ%��V"� �>����r%�bX����6��bX�'���Y��K�O�Ic\������9ı,O��~ֳY��hј�浭�"X�%��w�ӑ,K��߻�6��bX�'�뽻ND�,K�߻��"X�%� Ҭ�*�V%�J�m�HƏv��~���Uj��wk5��6C!  6�  pnۛ�����5��S�S����:&��V+	ح��l��y^s�تb�mk�Uc�YQ ӂ$�Gg[����N[���F8f�9�-ۖ�S.�x�ڎÎ^��.�y���t�qm�Xg�\�tF���ɱt��@�Y4��S�\j�!̸l�6d��;]�=����**�IѬI�U�bg�.C �ٖL�4��k.��S��7Dr���iy��K5uasZ�\�[��gs2�FkR]h�jK�h�{ı,O���ܳiȖ%�by�۴�Kı/~���r%�bX���xm9ı,N�5��5�-�k.�fӑ,K���w�i���S�"�j&�X�����m9ı,N����"X�%��~�,�r(~��DȖ'�Mv��u��f����r%�bX��{�[ND�,K�~��"X�%��~�,�r%�bX�{���9ı,O~>�d��j�rꙩ�sZ�r%�g�,������Kı?}�ܳiȖ%�by�۴�K���12&~�kiȖ%�b_O����F�&�j]�3Fӑ,K��w�m9ı,O=�{v��bX�%��w[ND�,K�~��"X�%������.�[V��u<���b
˷��n������a�4I�WFfh3F��(͛�a.����2L���i�Kı=�_�]�"X�%�{���ӑ,K��߻�iȖ%�bw߻�6��bX�'�5'{�a�֦j��L�֮ӑ,KĽ���i�U���Q���ijW b�ʁR�R '��W�D��L�bw�{�iȖ%�bw���m9ı,O=�{v��%�bX���y��kS,֍�35�m9ı,O}��6��bX�'}���iȖ?��=�_�]�"X�%�w����Kı=>;����-֋MIu�ND�,T,N��yfӑ,K���w�iȖ%�b^��u��K���ȟ}��ND�,K�f�g�al�]h�5����"X�%���nӑ,K��ﻭ�"X�%��w�ӑ,KĽ���m9ı,O���.wY����5���/ꞇ����ά�]Ga��,S;ۣ���-lD�͉	�c��{��7���}�m9ı,O}��6��bX�%�vkj'"X�%���nӑ,K����A_��*��U�M]�/�)!I
b{�����,K�߻5��Kı<�]��r%�bX��}�m9ı,K��>��ѭI���Fd�Ѵ�Kı/}��[ND�,K�u�ݧ"X�>�>	F�!X#;��a��df�eH�H��IH�"�`
@��RD�c	��hJRU����ů�o��|O�|=Ipc�l.7�k��m�z��z4("B�b�R���iY�%%B3瞑�F0�(J²��qS���!HЅeP�A 3ԍ#1�b@���@�"FP�aB�)�*��,R!= �4֘Ԅb�}�@j�F  �`p�]M�]!��D�*B���
5��������si��-�����y��(p�uZ�++����|\V��%!I$&:D��7���a!4F��d�3A�鳐<�F|Ah��p@��≡S@�T�PC��Lh(�Q4 iF�	"y�}��"X�%�����"X�%���>�Ma.����2Mk5���"X�~P dO~���iȖ%�b_���m9ı,O}��6��bX!b^��f���bY�7���[}�c���eh�����{��%��w[ND�,K�~��"X�%�{�ݚ�r%�bX�g��m9�7�����7����U�t7%�n�ؑ���:����xzط-du����V�w�{��2��je�ѣ1�f���"X�%��w�ӑ,K��w�m9ı,O3߻�ȢE?��5ı/�����r%�bX�������-֋MIu�ND�,K���Y��Kı<�~�m9ı,K߾�bX�'���N@S�"dK�f�f~�Y0��,3Yu�6��bX�'��fӑ,KĽ���iȖ%�by����Kı;���{�7���{���u�O~�����ͧ"X�*�B+�3�{�[ND�,K߻��ӑ,K��w�m9İ:#��D�dXi �(` jD���ͧ"X�%��|}�٘2�ͬ5�������ow������r%�bX"� �~����i�Kı=ϻ�6��bX�%��w[ND��7��;����{�����'P�.���r]��d]�{-�GgX���k���N��mv׏�{��B)9�t�s.�jIr\ɗ3F�ؖ%�bw��,�r%�bX�g�w6��bX�%��w[ND�,K�~��RB����b�t����
����2D�,K����Ӑ��DL��,K����ӑ,K�����iȖ%�b}���ND�,K�橫�L�%ԙnk6��bX�%��w[ND�,KϾ��"X� "~���fӑ,K��;�ٴ�Kı=���gndՙ����3Z�ӑ,K����iȖ%�bw߻�6��bX�'���ͧ"X��>����r%�bX���f^h��n�ZjK�h�r%�bX�{�yfӑ,K��>����Kı/~���r%�bX�}�xm9ı,O*�v���Y ���m��v��k�i�k��HH  9��� �0�sfq���0��-q�xsu�k]���ZH3�;Q�ѮN�Z���v�\.���u�D���ݢ<�헴�ol9�b,��L�`�hc<�EP��8獞kl�7qiڳ�]��B��;v/:�`,���Ti��p�m�7Jt��uӌ��c�Ō씁y[S��g����{ǻ��G���V׭=p�áz�J|􆣗�u�ǗN�ln��8֌�,��Bk��E9���s	d��D��e֬�v%�bX�Ͽfӑ,Kľ���iȖ%�by�����DȖ%�߻��m9ı,O~����3Z��5��W5�fӑ,Kľ���i� X�%���w�ӑ,K��߻�6��bX�'���ͧ"~A��2%��������I��5�������o���m9ı,O����iȖ%�by�}��r%�bX����m9ı,K��>��ѭI.K�d�Ѵ�K�� �w��m9ı,Os���ND�,K�߻��"X�%���w�ӑ,T����i���M��XUMUɐ��%�by�}��r%�bX���߻�[O"X�%��{��ӑ,K��߻�6���oq�������y`,�sΤ��i(;+Y����r�V,�IF.آ�H7m�띩���l[ ��w���oq�������Kı<����r%�bX�{�yf�9ı,O3߻�ND�,K��]�v�MY�ՙ�.kZ�r%�bX�{�xm9
&)?��J?�6ș�����ND�,K��fӑ,Kľ���iȟ�(dL�bz|~��y�3E�M��Z�r%�bX����fӑ,K��=����K�2&D�~��m9ı,O~��m9ı,K�Ӷ�	d��D��e֬�r%�d����"j'�����A'�kbH$��=�I�$���~�,�r%��{���u�O~���³�����Kľ���iȖ%�a� �C��ͧ�,K�����6��bX�'��{�ND�,K�;�u���ɭ�f[s$�t�)^e6�^�C�=���m��ǉy'"T�Ψ�G^�r���2�͠k�����{��7�����ӑ,K��߻�6��bX�'��{�_�
�"X�%��kiȖ%�b_O����F�$�.�3[ND�,K�~�,�r%�bX�g��m9ı,K�~�bX�'���m9�A2&D�>����]Iu�\ԙ�e�՛ND�,K�����r%�bX����m9� �S"dO}��6��bX�#�ߤ�_�RB���+�r�nʹ	�-�k6��bX��>����r%�bX�}��6��bX�'���Y��Kı<�{��r%�bX����3�2j˚�1��k[ND�,K�~��"X�%���߻��6�D�,K�����r%�bX����m9ı,ON�{�+�4�k�ݧ^Zx����'�����sĦ�u-c�N�VN��J帛�nŭND�,K�~�,�r%�bX�g��m9ı,K�~�y"X�'�w��"X�%�{�~��Ɇ�VZf��Vm9ı,O3��6��bX�%��w[ND�,K�~��"X�%���w�m9�@$ș���~���1*�L#?=ߛ�oq�������"X�%���w�ӑ,K��߻�6��bX�'��{�ND�,K���Rt�Գ2��չ�m9İ�Ir'�w��ӑ,K�����6��bX�'��{�ND�,�`�$VAB
��dK�~�bX�%���gr�֤�%̙s4m9ı,O����iȖ%�b�Xb������yı,K����ӑ,K��߻�iȖ%�b_'��K���۩�Թ5��'m�nu�X���`N8�m����/ڢ;]nK�`�\[����{��7��<����r%�bX����m9ı,O���6���1
y"X�'~��Y��Kı;�ԟ�f��֦j�u%��fӑ,Kľ���iȖ%�b{����Kı>���ͧ"X�%��{��ӑ?���A`T5Q,N�~.�?�d՗5.cL�k[ND�,K����iȖ%�bw߻�6��bX�'��{�ND�,K�ﻭ�"X�%�����^h��u�IMIu�ND�,O�� @"~����iȖ%�b{�~��ND�,K�ﻭ�"X�%��w�ӑ,KĽ����K&�Yi�˭Y��Kı<�{��r%�bX�`�$�~�ki�Kı>���m9ı,N��yfӑ,K��{��������5UT��)p�[e.G� ��  ��E��٥t��p��S���SA�zw�I��� V�pg�em��˦;wD�b��9��v�sPlY���a��������#��c:�ۤ���t�n���38�c�mɹ���`���/��8M���-�x	����V�%��-��8%MF5v0���Egn;=n�x���n�O��\�ש��p�n}�	e��<j�N��5�rn9�}�ݵ)눕g����%�bX��{�[ND�,K�~��"X�%��~�,د����ACșı=Ͽ~ͧ"X�%��t�����K3.��MK��ӑ,K��߻�iȖ%�bw߻�6��bX�'��{�ND�,K�ﻭ�"*~!("X���w?eѭI.K�d�Ѵ�Kı?}�ܳiȖ%�by�����Kı/~���r%�bX���xm9ı,K���t���Z��3$˙�6��bY�*�@� ��,�E"���o��ٴ�Kı/�����r%�bX���xm9İ?�	�?}��Y��Kı;�ԟ�f��ֲ�Iu%��fӑ,KĽ���iȖ%�`	� H~���6�D�,K����6��bX�'��{�ND�,��w���~�x˩VլV�n�-�md�%��V���a7m��#ٮp����y	4[�K��2�Z�r%�bX���xm9ı,N��yfӑ,K��=�sb��E  	�L�bX��{�[ND�,K��ٗ�34]h�u	u�ND�,K���Y��>G"DdD@8�iș��>�Kı/{��iȖ%�b{����Kı/~'m��f���e֬�r%�bX�g��m9ı,K߾�c��#(.�j'߿p�r%�bX�����6��bX�'�Mw2�.���5����Zͧ"X�%�{���ӑ,K����iȖ%�bw߻�6��bX'�`1"��=�~ͧ"X�{������;�V2��e�����7��b{����Kı;���ND�,K���ͧ"X�%�{���ӑ,C{��;���L��ʶk��A���db�ٮր[���˞,I�T��Tןw��w��;��j��eѭI.[�&fh�yı,O�w�,�r%�bX�g{��r%�bX��}�m9ı,O���6��bX�!��w��ła�Nȱ�{�7���{��g{��r(���9"X��{�[ND�,K���ND�,K���Y����oq�߿z�����Kl[ ��w"X�%�{���ӑ,K����iȖ?h�H�c0�*[XāH� E��� 6���hZ��I�2Y*��!%c IZ�DQ� �#�<�����ND�,K�����r%�bX���ݽ�5m֥�e�u�m9ı,O���6��bX�'}���iȖ%�by��siȖ%�b^��u��Kı<=;����.�h���kFӑ,K��w�m9ı,O�Au����yı,K�����"X�%���w�ӑ,K����w/2kZֵ��3WW7�l�=�p\cMՄ�3l�n�um��zqQl�B{=1��(�=ߛ�oq���3��m9ı,K߾�bX�'�}�@AI|��,K����6���{��7������p�V�a�����bX�%��w[ND�,K���"X�%���w�m9ı,O3��m9 O�W"dK���)?Z�fk3Z�2浴�Kı;����Kı>���ͧ"X�%��w�ͧ"X�%�}���ӑ,KĿ���]�%̹�ff��"X� _�(�'����ͧ"X�%��fӑ,Kľ���iȖ%����",`�!�R'{�8m9ı,K�i��u-�j扬�.f��r%�bX�g{��r%�bX$Ͽw���D�,K���ND�,K�~�,�r%�bX�����r�˩V�k=�ZM�	���M��c�FꜩF���v��\����E%���ۚͧ"X�%�}���ӑ,K����iȖ%�b}���ND�,K��{�ND�,K�O��ܳV�j\�Y3Z�ӑ,K����i�'�@ș�����6��bX�'�����r%�bX����m9ı,ON�2�Ff��)�u�Ѵ�Kı>���ͧ"X�%��w�ͧ"X?�.Dȗ�����"X�%�����"X�%�~����ZL5���5�Z�iȖ%���"{�߿fӑ,KĿ~��m9ı,O���6��bX�ȝ����i��7���{����)���k����̖%�b_{�u��Kİ�U=�xm<�bX�'~��Y��Kı<�����Kı>]�`A�E�@ ߋ
$O�#�� i$4"�
2�$H!�$B�"E EK��F"0 ��y�LM�`� ��{р@v��#
�T�$P�k
��[BVP�!@�X���cWj>"bF$c�HD���f(�6J[p�B! qq��$Q@��@� �b�"A� �X�륕\c�F�v<*���𜊾$�P��Y ��	D$�#ŅBHń$H��$�0Hd	H$�H$cRT���kZր�`       H�%�i.KNkY'4l0x=�@T�'2<�@At��'f�i�f�        H            �e�             ���  N 8   ��p�6�4�$u�s�N�z���}�Ӫ��I$�)��c�9�:�#F���ۣto4ȎìMm����Yܓ;vù�@��n.�[9��������t�m��8뱟�[n��e'��n��zc7I��:�wnc�>�)�÷bGW`]G�*���;t���v֛t�%�,�x9�lv����Hi]�z���x��\�%)Πs˧������S�ciЌq�D�Yx'6VZ�16��j�=clc1:!�����v�vθy�v��n��\"�:7g�u�&�k�&ݲ�<�t'�ו�9�{u��[<b�ZrN�ecBd<�N\t���x8�Η�s����C�m���4Ѱ�nj�����=��mg������S��"j�y��v���� �ٳ�eo@Ok����K-#�ܞ�f���c��ҡ�3ñ�L�u�Q�vp07�t�� bFҤ�"�4�R�k%����)�d[��k�#��6l�]Y�s����v�z�k���[��p�8Nw^�*����Z٥Y��={6|�n��:I$�P;m�Z�k�NP.vPڪ��	��[7u����at�h�ڱ	�Lp��%[�t"��r�Y��S:����󲆇Ɨ��跶�V�4�S�Wz�{k4䷧N�;N�$����a�l�ڴ�d�Zg��fh����]��Wd	^ h�����o<uu��vp��Z�"^�u �`P���:�a���;��t��IbԲ4v�x��X�8��Z�%W����LOs�4��M���#˹��������Ns�7�P< ]5��p��X�(u��Kf�Zԙ3Z���TeG� z����
��W�� �	 � �ډ��
*/�_5��kZֵ�k[��iM9��ր��� m�  ��
aa��ݧn��t�g������Z��(vvA�J�<�9mǒ;m��9����I��Ǜx����ŝk�%V���u�T�m�^�V�tg��8��ռ��hc�Obzm�:<�kd�T�/��C�'6�Gٹ�����nSj�Rdm֜��;��.�;����s�k�R��ҭ�Tk���K���X�K���;9�g�[���65��%ӎ���Z�\�]h����SȖ%�bw��iȖ%�b}���ND�,K��{����"X�%��kiȖ%�b^�S��.�jj\�\�33Fӑ,K��߻�6��bX�'���6��bX�%��w[ND�,K���"*�G"dK������n�W4Md�s5fӑ,K��?~��ND�,K�߻��"X�%���w�ӑ,K��߻�6��#�#�#�v0���(F�
Iǿ��,K?
��:���~��ӑ,K������"X�%���w�m9ı,O3��m9ı,N�>7or�[u�sd�k[ND�,K���"X�%���w�m9ı,O3��6��bX�����M���.Z���G$�A�q�����L:��NK�\-����/m���S����{�n8޹�LNAG&x���@�u��=e����T��Xnvo3Z�՛�r��ٿ�����F�)�P�"�S$1��h�&��C5XB6��I~���tD|�����x��ذ��F����\n17&GR= ����^,:/�Q����&��}X�Sk���I����={�Q�x�נ޳@=�Vs�L��q���Z�7��L�/����ﾯ ?���=��d$m�HD�Iv^;Wb÷�����>z�!h��\/rk�q�:��a 4�F���@=�f��u��Q�
^���d�R��+�.���jf�� <��(S'��X��&��@�vD�DIH&��@��'�{��ܪ�!��R�DC=j�&��0uGJ��_%
?����~�oՀﾼ�SuYV�mMYjU�uv�?�DB��ߤ�=:�����I�%Z��, ����ԦQ�ټ7�w!��� �^`}%x����h��fW��6�$�<�p��6�����ƹ�Q�'Sb�7��Z޹ڭE�4���bN)�Dӏ���hw]���$�D(�D$��=�V ��(�d�W�����W��Z).��k���D�b kR|v���.�jj\�6��������<]���@���=�56L�V�����0:!B��P�o��������Ł��$�(���F�� �u�R&�bCĜ�@/u��W�%z0>R]`��fg�#�<��Uf��	9�������va�A�&�fݖ2�y�c��'�����������	���I8���nh��4Z��Y�y����cS�ŐQɚ��侈BQF��}X�w׀n�ŀQR����c�����z{��=���m~���8�uu��	)�o� m�, �-נz�+XP����nM����^Q�~��`�w�LF�Q)C�$#��E!(�D��q�����@�UUO=���2 뮗!      �n����/;vH��٬H��wk�-���VNy�;sۃ�=n��5kS`ګ95��/k�r�J���[�m�"�,ڢɍ������]ڎ�'p�tWk������۞K��b(G�I�&^�/;��l���G�7B֑Me9��ϭ�ݷ65mv��;.m�l@"pS�:!�:�[G�� ��?0�	 �HHAP � �D���t�:�,�K�k�<��;\��qx�α�����n���&��n���N�.��л+-��(�?Kn����	~�m�,��O�DFG0�n3@�[^���f)o� m�, ��ӕse��$v$���Y/0$��>��+/#��[^��vA$4���p>���.��,�vQ�zu�����o� �k��*�M��-J�n�� �^Q�|�F�w? >��wu��;�߫`���	�Bn����zCtO>���.�ֲ�;r�=���k��x�&9�$��<Vנ�����{��@�[_�jbN)���Y�$��~��TS*�tY��͚����<]k�=]��(L�n
L������,��ge�V s�M �=Yε2C"r&��3@��X��Ku�Y/0=%x���и�%Ⱥ�]�UUр?Ss�t$��}���s@��Y�g�ܖO�$��&<�u���앣ƍ��ۡ�ۊ��y��n73s�2(F�bD������h��h��4�h��*��$��7w�=׋9D/�EQ�w�F󯾜 ��hg�սs��&,��L�/w�ɹ'�g�]ϑ�"M��0	r#�BH�gw� ��ŀP�]"B����V]�BP�{o�p����ŁТ"'���`euT�UM����������� �"�o�/�s}�`��@��_�>d�����~R6�ňɵ��˹��m=�u N뱝w�MŤ�W��qmY��M��[��{��@/�� ��h�V�S$2'#@���^�g�BK�(J�>}x�w׀=׋ ���.(���a 6�f�_m�{]�ВP��7ذo���C��\�۹�,����y��J�d�G&���I0�0P���?g�_:h�r
�D��7�CRM�7� �
7ߨ���x �]�����UG*ڷCvn A��O����ƭ���ӃHt�����PqnxVnHͮ9�5v��� ��� {����Hn�fh�������0L�H� ��f��G�BI*�������X�yF���_�jbMƉnM ��h�n�{��@=�٠{��U��91I�SUw�В����~X7�F {�� ^�4�v)���6�h����}�(�����w׀{��ͷ��@�UUO>��qm���		     �)�^�FعfΖ^���GdL�(��6�D�:ݫm��:p�l�K�z�l��.:wm��`@*$6��\��6��諪�"��g)�7l��c�
^[��O	�͑��f���l�J������$�u�/` Ԧ�g�#`!�ʼ]tб�鷵�mv+�=�-bt�m��u��c�9�lel��4��@Y�:y�7Q�֨ssd�Y��pϷ�Ӝ�՛�ٽ�Z�4ݫeY�6���y�Y/0=�^0,������_�u5�j�tIsZܓ��f�(!�T\���b�>��(�y��<֫%�3wrUA53wX��,��2n�^��y��V��j!�b�D���ߡ(S���0w��;��y�X�ʕz&DL�Ȥ��}�h߾v����4�u���9��l�#^�/m�cvYyۢ3�!��W\��v��\��b-�a�����F�k��s�h��$���V������>_��׀j���u�˚�u����nI�>�f�<�����w�(�{]�w]g��)�i�}���Лs4��Y�{�hwW�y�]�����J!I�@m���K�Uk� �{��������h�=�I27�	L�hwV��Ҽ`Y+р}�y�e�)�q�U�kڝؖ��C���ن&��,�7�Ю�y+��5�o���xz�AW�[�����^��K�
����{-{Ģ&,dNL�/u�h�����X�kŝ	%
d�˦z��.KRdNFh�~�]��٘��33<O�
+���	$Y"�<.�W�f���$Y��b�i��K0(S �H�n&*�PR��Q"�@�>^��i��9�`���$�`B���¤��)
�J�����(zA.�!)�F��&*B���	���kw9c9�0������)�7x����ڍ'9�jF!���2X��1��ʇ�D��2x��ԇ�(JF����,c2�c
��+(J�h��|�06�Q���� 4�@d"*��D}D=@4�&�F
)� �_�؆���j��DT������0̭�_�70mƉ�M���=빠^ה`r��
g��x�jzWU�tUڛ�F���=�^0,���>����K����C��m�9Ȟ(D�`�P�M�u�.u�Տ�/���9&*m��/k��zlW��Лs<�~�h��4
�������������O�D�B��6�f�~�w��'��N���^Q�j���d�y��NM����n�ى(�o�$��� k��Ӫ.f�䪂n�p6�`�����(J��UF�����rO='�]�4[�3Z��]���7[�0P�%������ ��s@���V��I$c�bs�sы]���7&����.�I���pv���ې��2@L�ȍ �hWj�=��h��4�����6�D�G&���:DL��ذ��L �n��QVW��&,�@�۹�w[���
��u��� ��Fӹ�v+���$���В_D(U��ޓ ;����ڴm�����(%��&7����B�_t�_v,u�� 6 F � .��@#3���>�U,E%���UR8�� �� 8�/]є�K��^l�j���uH�h�Mʍ�f�7<�N�Z��Dun�u\ct�l�S�xi%1<[�k�+\�Y����lMnx�a�r�:���wmk��L�&�L�z��J7-�wl���&7<�K3�ۅ���M�,��!�J����Lur�tO�w���ǿ>~w��u*ѭa����IP;c[$�5�:�u�s[e���:uv~����'�|�:�I��\�λ� ��� �o$�#􁯺��Ϣ6D����ԉŠ{��h��0���^�ϔ(�=��3rUܒ�����wwd��n�/]`�w4r�J�"&L��#��[0/]`��`tB�����`�uT�����$j94
�W�{��hۨ�z٠{��x�;ndM�'/����u��ٹA�p�&��X��M��2C����#&I�mǠ{��hۨ�kw�K�J?�
6����� �t�����خj��Xm���pB��			"�Q
�u�xO>���,��B�Q
LR`�q�[4/]a���%T��`}��&�Hn�s����W��=�w4m�h�l�:�dl�I17�m)��o�	%�I/���I��}x����r�=rI$�A!�nL %�ڸ}x�sŋ���7�8	�4S��n�SpFi�4m�h�l�*�_��ٞ �~��;>ϒ��2d�������ДB����V��,��L�m~����$j94
�W�{�w4"WKm��M��j�W755e��EU]`tD$�u����� �@��z���u��G$Cf�c�Z{mL
�����x�����;����Yu*ڴ���9�a�;xѝ������!ets���to���������&7�_���*�^��w4m�h�;�29�BɌR,��X�kŀ6�I�~�k��J$��\�SM���x6��@��ۚ��0>�ʘYu��aj}��r7zfU5v�>�J{��I�{i��^��z�_F���V(7A�Aˀc��8!�!�Mb�A��I/�$��� ��̺�h�-Z�4]�ܘ�V��>�	%�ϫ��ذ���6�������*���z���K��Q���;5�×��O۷1���Sv�*u�v�	!$�@��z����-�Q������-���ϤJ6��&1���qg�'wvI�{i��^��IL���'�i�By ��F����?��䪽^��}���?��PLRb���0>I$��m��<���o �x���ő�B�ZW��?y�Xm��Z� �
�A�	�����U�������Q�
�� �l  :�8,�s&\�*r�';#���(��6m���ZS�m �*�-d@��X�
u�3"�k��7^��(3�˶�%�v�,�9���ш2���a�0�8�\��k� �v�:l��ݍ�R��a!gU¹�RG#��H����Tf.泖h�x���^�s�ڬ[3�(۳�zqQ�媪ͺ�S��ĩr9��s�:-]�֔ӋnmqOWa?{�����>�p�n�ݰ��0-����l��U�X���c��Cq%��I���4{eL
����ּ`{.T��i���jh���0z�� ��>IBK舅Z����}�`emT�UV�j�.˻���(IOW>��� �y&���@�ve�(ڊd���z����%
;��I���p/]`����'R��K�k�2E�	��<!�8����=�F6��pn�뎼O'L�ѱLi�[kC{eLz^`}ex��J[�0�u��D˙�7$����V�
��K�$�����7��`�x��A�dq%"�b�h{�hY^0>��0'�T���Zպ�]v��Wx�)�>��wvI�o������=�V�1(���2G&h[Z�*`���+����Wa�[^"n��g����{ss��ty4�u���v������� �9�]uũ��7ծp}���^/�I%�D(����&��S*�A5ee����\�<�w4-���}V�$T\>Y�lQL�jI�}~�s@�ۨї3��D0(�M `�� &(D
��)T]
����g�����������Yδ�D
G9��ֆ�j`���^0%���\�KUv��5W& ������/�!_�������� ���0�J!D��Nxx`,�s�f<�i�4G�0t��n��n+N��5�[��nr4sF�Й� Y��}z���6T���u4ڂ�b�ɠ_l���3��ď{�$�9���������U��ӗV��N	cnj4Ϫ����/�S@��*U��&L��#���8��x�`~JP�BP��PD)���I�|�꩏�U���EZ��� �^`_^��+C͕0&+w�]|U�vK���ITmv{�8nLv���S��]��[�FM�F���=����.�V������0>��0,�S �^`=Yδ�D
GHh^�������/�S@���q)�E1G�MUɀ=�s����{z��=ϲM��׎4F�C�C��C}���?���4/]F�y�Z�e��j
I�<)&�岚���@�}V�=�ߵ�&���|>)b�*��0!������2��݄<���G"�!������ ���ENA���"J�KebB����%v�`E���6��(c	$aG@#�%@#��*8&����6����ٱH)���!Rdl�����>���S�Jw���/��   $       A6	����ɮ��Bp�y;�0
�%�5��V�36m�      ��            8$              -�K�  8�  [2+����mպ1��]��ݪ��os�3�N�`3"S4-$W8z�uv�N$�l����{c�;�	�rNn�Vg�u��n|���Y-�s^��5��D-�YIy�ƌYu��4h��[�g���{f�F��Y� �;m�3��m]����UR6�;�U*��C�MX��`,g� ճ�{]=Vmv<�)�-s�'���k�ݝ���v�5�d�LUK���Kۯ6��g-c ���ѵ�2��S�UK;^k�ˑNJmo�O�{/\򲑬�E\�����f�ݷ6˳�T�v�ځ46��ݳ�L�q�ݸ��;qև�خ���v�`{ۍ���c�����6ٯV �{;sK�@(j1�]�����`֢5�T�<�pݣ,�F띘ݮ���훨m�7lp�v��t`&ص��]�*�wm��E��9���^A_%p���@���p�Yt��7&�qҐ����r��a@��-�&�뭧uЗVS!u��rt�Oh��<peӶzy��n� 6�4���蓮�צ�v:s�
�>8*���-Tmk<-���uz�ڪ��������S�S�Q��#���ѻ@J�TPN+ %DW;cRq�Y��ݸ���n�i�
����7'b;��9�xKs��+�Z8v���`�'���k����р�gM��Q�c�[�����od8��h4 �iQv�!��m���5��Ӹk���,���{.;,'O��l<Ld�gT
���$f�n�fW�^����ZU��*��c�8�o:6ܦ�']�!W����m��3:�\�;�䗣���w=�cnp�ݔIQ���ww���w5>OGh��]���q�����{��|���UU<��ln[V��\�� �  p!�/]Y\vĺ�U����y[�]$��zq�k��G��<g���V�m�k��nP����t7g�-f,��8�p�q�Cs���Nh�	#7���%�8*����@�@����f5�8:�w[e)��lk�V�f�[��+��6qؼ�4c�r+Z��-�tMgAs>h�
sG2�L�5���M[��1�Jո���1n�[�m��\�������ژ�ǂjG1(���0m��=�uM�0	%����eJ�oa�����CM�0	%��׌��&tDB����9UZ	�TU����o�0>��`}�^�	6T��&e���)�cn94-�����hϪ�{���Vs�9�	H���0>��F�j`���׌������S���f���b<g�[4����(���)�ڰC�d�v�g�Vj�)^}ֻX+�t���<u}���]�m��(P��u�Y�}���)1F��E���kp��)Ŋ�P(��FF+�E�����B`�P"�<� �Ui,�}���:��h�տ�GԹ���PRDF	��	���������mLޗ��V�1(����ɚ��Y�w;g =�w����� kWL�Z�V���6\��ηX��S}����b�?w]f�ؽG5Y#m��	�S�Y��0[�l݌t	LW�����V�v|sI��nڔ��`.��{7���{���׌��F.�����,�lQL�jI�{[Ŝ����(����{]����Zs"p&L��y�u�.��ُ�X�D��$-ߦ���}��u��S)��Ӻ09DB�O��u��[ŁВP���![��� �I���t��7T�]L�� �����`}%z0*�� �o}��R��+�;�J�m��ӳ,Jn�g	��`�.�uUU�g�E,Ti�Drh���<�������<A��wa��d�Q	�/͎L�/u�o��(Jd�}Հt�Հ=o�әyx��$�a���*�^�Wuz}���<���9��0ⶪa��A7j��WwX��	W���`w��=ה`dBJ&�B�z������<��{O�آ�&1��z�h��4
�נ�� �=��v6�##"x� �dbs��tX��n�j���;��;��պ�˞���Ɯȅ	���}o������w����w��>���3tv]"�ս��n�%�����W��؎�c�<Q��hiH��Y�=v�9)�o����V �m55Sb����/YM���*�^��Q	%3����wN]�3rMY3EU���FR�`������;�� F0�#�
��1`I�d�B��!U@ @���H��D B@��@ ����2B �@�$B	@?�?+����v��Ɇ�.����   ��kM<�.��q��.��9�5���F��Dχ�t�;a�#m��i��Zn��[�#	��V�;��8�v�\�=sjt�-���9nZ�D���It)����d�.s���c��`޺Sw����ۄ7�
ӝ�<ٗ-t6x�7ܗ �ΕK�M�ь�55֜�5���k30���GB��s�*��s7���=�n���Ͷ���r��̓���׶u̿��s���gC��.v����=�y�e�0>�������&1�rG���h����u��n����ɲ4t��.���I��$�>�O�����1/��������c����Hht�FR�`�������q.Ў(��ӌ�*�^���]���_�Ɓ�u��nPL�nDB!��/��%՗lkl���\unq$�O\�7<7;3�mH��o$R= �޳@�e4=��*�^���p��j
0p��krO��_M���DX5XG"`�1aB!
Zߟ M�v 8��B� �����=�w�n���^�{�Y�{���	D'�6UY�~��� s���L��� ��Ɓ��J����	�ȍ����/0,���J���6n�����v��Uuu��w�|�{�/�y��0
���;=|��v6�2L��Bd��#��u��5�ܢ��2p;v�kr����b����:�5�1��������*�@=�@;=Y�1̈Q�b�Nf��u���X��x�x��%2oT_�(�8��<�F����Y��5	��� �EF��lYJaB��D(�i];o��I�j��X��#o#N=����b]o�@�<`}%h`U%��[�F���V$�� ��,�o�I������4��|��q�$��q�%]��M����c�m\=<κ7�/�݄�i'�693�=��F�Wuz�u�J���ذ��=��˔]�2YuWr`w]g�BQ�Wa��X?�ŀ~ށ ���8��Lc��@?��`_Z�����T�XD¬���(�I����/��hw]F�Wuz�6�:\P(�~�krI��Ͽ�ȅ$Ɋ!9���Q�U�^�{�f�}�s@��v�&70�"�t���4�^�4gn�H6<���SXy�{q��v���I�F��M�hwW��^`_Z�����1���n���
��� ���2v�b�<�d����n[���PQ���������+C�.�Iy����>�jKxK�����J���K��^`_m��=�*Wf,��H$B7"4
���Iy�}k��V�R%s{��;:�%��Zl��  v�  X`�����I��l�ej;;���[L'mp,�ӊ�s��M3���x�]&:7L��]�s��yWqIu�;v���n��Ey�0�o]#ND-����o�=y�γ�+�V㈝�SkQP7q��
��1��X�N.��GK�:׹Ʊ�d3[�u/�C�����j��.X�w}�ww��/|]�~J����\<3�F�dSҝu��HM���9۷Q�l�p�ؕ\u��q\��g������}k��V�R]`y
��lx(�I����/��hw]F�Wuz�f�vz��c���1D'3@�Ҵ0*�� �������q(�8��0i������z��n��ub8�������{����zV�R]`}�G���UVm��p���9�xwHpNεv�[N��K�k�z:��ݡ�;6���`_^��J���K�ޗ�{
F�I8%������u��~�DE�����DHT����� ~wM�3?~H��%��Y!��$�����`�����Fޕ��}�tYA�����1��{�Y�_l���u]�����Y�<s$�ڒh�ـtG���?��� =�w�t$�}����'R��K�f���t�v�ɔ�a�;��ڎ�n��pkp�:7OT���]r�.��=/�C�n�z^`Yz���\J0�%0i���������ـ~���:)���v�d���#����/YM77?bm�ѡ�c]�{�R6�s�]�IM`.(8���@�ZC���#B/�������*��
�
,j J2�eŅaF��L(�Ä��<����d A� <C3/<cqap�/�x' �o�
M���<�m�R$]���U���(@�D$� ����1�`G ZƄ�@�h��)(���*��B*>�� ��v�p"��>P](�� �����/��*��P��Q<QH`:@��Q�r�@��ji�8	�0,�Fޕ��T�X�/0=�)�F�y������u]k����f����puHM]�VG�t��F�˦w^�8�#�m�ܚe�2�ڳ��t�r�s�\\un�`������>���
�����Ҵ0/�n�(n����9�H�
���/YM��Q�Uֽ�qW�1ǂ�d���z�(�����T�XIu�L�%�7�bR8���4�]F�WZ��Y�*"/(�/�{jS7Aus6ASUr`u��:DD�}���� ��Q�RÄ�;Pr	��$��&���n�8;9]�ݦ�+�<���ަ�sV���d���#��f�z�h޺����ܷM6��&���l�J&N��&��� ��C�Q�<��I�@���hu�@/u��)�{r�vb�$"#�7`U-�d����zSX�͋(7���9#��f�z�h}��ηX��!!B���8�P��r����kZֵ�W5�ˤ�:�.B@   �v������C�;��m\��竗p���k�E��:NE^�7�^�5Lmzv�����c�������a�pNf�[lu�9ݺ�N�Ӵ�\����v����j���:!�-��s�C$��������c42i�����a��R)���x��-��5�uڻ&'	ڳ�H{*�4k^(�AT�N��|�d��3$̑#^�N�����N���WR\�ݒ2n�W K��#�G2)�nO@��|h{�z]k��f���9׉̘��b]��
��XIu�Y/0/�S@���q(�8���"z]������zU�	��o�y-2c`�q��f�}��^�O@���ۖᩦ�`�$ӓ@��F^�k�.�-��v�7tB��!�ӣmN�sz�5�'n.��l�b�q�L$i�F�Lvy�m2N�zm�m��\� �u� =n�P��޾0r��R��U�3t�������J�BV�b�P�J0�� {��ϵ�gB��Q�%|J�j�*�]]`��׀?;f(Jg�_M`-�`�\�;��uj��wx�OogN����נ��g�9׉̘��bQ�C@�ҭ`U%�e����F⩧g���ç�ռg�[T����Q�/�{p]v�����:���t�ζ�2ԍ&�
���,��ר��ҭ`LFu�ƜI�1�i8���~���bG���ӯ��;���I)�yw#&��l���&f���޾0>�5�J�(P�!�"��6f��}�܁}�4=u��"?D�p����ħ�_M`-�`���P����߳�ً$0�$��'�*�@/7x�`}�k 䒈�[#��.�\�ŵ�.�����n���&a�WFڸ��q���e��;R㭗�3a.j6����^ ���k��Q�K}X��/�L��a&1I4�ߒ>]~O@�[�����ל���LJFLQ�0*��XIu�Yo0/�Q��?��JaJ`�=������?;f�(Q	ZQN��k ��ZݘӉ����@/[4��*��z]��[r���6܈��W;Qv�&�(X�2��3���7H��]0FF��mD��iɠ_l��W�S�*�@/[4=���"?D��zU�
���,��ר���Evb�B"<�q=�����@��M�z��__6,��LC��ګ�� z���ـ9����?;~z"����Lb�h�(��ҭ`U%�e����������1x��t�\�� �  p����՘F���S��T���Gh�ƥ]l����9Nͣf <���P	W=��8���:x��ʵ;{z�r�Zs��[��C�;���1�rr�P�Ӱ2u�Γ�WR�G��d��;U���^�U��)��gFJ����;7n:N�(X֬�[i�)s�h�s�{����Ȼ<4�iӴ���<B�L=qv���\�������}�Y�^�L��b t�����
c��ͷ����Z��K��y�}z�����q(��D�
������e4
�ꞁ،�cMF�LPN= ��`_^��J��T�X�njmD��nM���*��z]k����p��ncCȏ�4�4
�*�R]`[���`\�J��*��s:��y]��&-qv6��2�]g��<�=��mI�ΐ���u�L��r� �[� z��]��B�!ӯ������y15jc�= �lۏ?f|(�,R1` mj��F������Q�T�k�.�<�R�{��0�����h{�=>���/�����M��sX'���C�`E�V�*�� ���^�뿭ģ�#$��u�@=�����/z�����h$m�h��}5e��*AV�:�g�˪㑠yglF�9#Ě����4�z�h�w4^�N���=�n�mD����`zN���M`U-������L��]7�V�JW$\����7_b�>���nz��2
��Aj	g�|�����p��1c�9��RL��u��w�=o(Jw{�,����d��I��@=�٠^�s@��w4
�נy�����m�d�su�/���t�5��{`�{l+=��sٸ�b&�� �8�G&�z���m��*�^�{�@�����LJFL\����k�R�`����׌+���#���Nf�WZ��[�:!%
g�v,w��E���J���Ի��{���^0=�^0� �}�C���Ey��~z���E�&�dĄ��/[����x��[�޷�H�Z�����0n:�d�cu=5�#:�qv�mtn�� Z,Y��&z7�
�o���x��[�޷�Z������d� L�"�f�WZ��m��w4}�s@��u0o&H�j8��}o0,��޵��n�<�T�^�Ps	1���/[��{�]k��J&w{� i�uԦ�Z����ܕV���Ku�{���^0=�~�����#�$�mi4&1�&�H�Y$���u1P�!56lP�+	R�)�HU��T���4LDK�%�4D�daHCf�0���x!Q^
��H�V凄(BHiS@�(�m��CJyZB0�!	YY`��ma�@���ӽ{�}��{���'��� �        ˯KН�Q2f����5��{E�6yU�l��{v9��hZ�      8 �             H              [��   H�   ��!Ӧ�����8Z�]���{�����;k!�6��g,�nn^u�����h��AR��u6����Y�I�f8�:�\�F/d�� 3l�v��*W;�]%���oLˣpT��1OS�eЙ�#��@zcY6,cn]:��.\�
�؞�a><����U�X�u������0R�c��s���a5��<\	]m[�ٌ�-��)�$n�,����A�ը�;j]����q�"�
.�"�f�v�k��nB^���6�g��`��n��EØ;b����pW��i��e�l����\i���Z�iӭЮKv�y���e��J.K����N��>h^k׭Kv�������a�֛����Q��xMM�N�ٝ�-q�*l�$=:1L���t6����l�鶷Vf
��s�M�9Áw��𜵅ua���9�cN���1݃6�G*�T���f���3�G�:r�B�Ɏ�7OC�����lmX���N���	ڴ���V�^��c��j�F�� Y6�`�C�V��j��uP;q/��b�f��S
etUVմF�{z"�ې�ð�B�dL,٢�m�'SQg)B㜱�.�UU�J��m�P�ˬ�is��q�����]�;�����D�c��x뫤�U[[Y���W�\�W,[U\7�v�*�T��r�n�n�����Zz�Փ����KX�ѷ2�dN��\)9���O��C�|��8�vӸ�l�K�R�1͋iSt�L��v]��D�r;an�B�(vm��V��9�!q�
�<?>>�s՝�Ur�8�����<s�H�]��.Y��i��#�]S�rs��]eSN�=�������V�W5��E��Q( ���¨Q8*tA}aP 1@OS�������ww�C�5UT��#$FI��	[@ �` �
u�وВd�E�nڷJi{�Е�1��Nf,ī<hzQ:��u�l�u�Kq�ێ:�-�O']�^6�嶈�ݫSU�%��lv�4���Vpvy�g{u�����l�gkb�̮�١ф�n<n��K�[���`���p�[Nj�n�l\�X]ͻan=�F����;G���Ӽ��(|#�U��<�S55�Z�34Mjh��6zr-V����۵��c˶�8u�̚��z����I�F�#ә�|��z���^0=�^0&#=on%�v��j]��>����׌zW�
�������M`��Iɠ^�s@�޻�]k�=�h��+sD~�wcޕ��n��o0,���p��1c�L�2<�ɚ]k�?�!$�Ϻ�ϻ�׋ �ڇT
iʶ���\<��+��'�:�,;�p��
�6��u�����m�u�k"L�Ͷ���w�=o�׋�BK�K��>������rh۹�?f${�w4
�W�u�~���r���2bn8���{�����'����`y��\J0��4�������������>��R-}t�jn�8a���=o0%���W��W�{�XT�$�A�"s"F(�݈s+��;Gn1r����{h�#��yλ{:jذ�`�5%��	ex����+.��٠y���D8%�,jL�=�u`/]`���5�Ŝ�%2{P�jvbs	0�B7&h}~z��4Y�(@�Q����L����HDd�H�B!��,��A"�ƨK�<�b�7��`�%����]��v�v�	�y�,���`Ee���� �7"nM�]��Д(�}�~�>� �7x�7�SstR��K�f�M�d��3�5�;�liݫ����&�v�5��۵�&��,�U[�m��ex��ˬz�`K+��K�v�pD����h�W��@��s@����=�g�cĚ��0bq�����W�Y^0"���r����IosY^0=ex��˛����"	���2TF!�Шh3>��krO='�W[���豩3@����9^�@;�f�׮�ގ�+@��(OВ`����ëx絤�7��d�f]�;j��)ӹ��{E�F����ܙ�r�^�w���]���s@�X�0L�71Lj9#`��Y^0=ex��ˬ�*_�9��ȇ�@��s@������2�V =�W�m:���*��M�w{��`yIu�O[���s���#�&F73@�wW��w�~��`z�`�`���P�w����6� ݤ�;9Qf��!  &�  ���f��nĕ9W�,���k����l��h�r<����]q�a��OM�f��˴�,��w=����A�U^{*��u�B����:U��]�����:�7<�F����u�63l"m���Ҍ�V���ASY58�]����4�ٝ&���r��N���d}�0�ۚ����w�o/f����Or���5ś����n�v7sv�<��+ѹ�u�m`Izػ8j������,�^/�D~��o� �܋�껒��&�ff����,�P�bG}~��9[���٠y�J�s"7��r����R]`���s@��:��bs	�&(F����k 7���[Ł��y��n�/�&L���qǠr�נ}���_��<��nh���b�����[l�/A�nq@p���g�v�W285�۝7u(sn2��1̌NF88ܞ��4�w4WZ�
�����h�&G��hܓ�}�f��D��j�K<�k�:٠{��hu��J2'L�UZ�=:�`|�a�I(��݋ �߷4���A&�y��z^۬K^0,���[�	���]�EMHM��5u�{[ŀr�o�/�l��U�@�+�F؄�m�HA9���T��t�d���ni;ny1q�s���y+�d�.{N'2'�ɚ��z^��z���p�ى�&L����R�`U�u��k���ٟ�"s��2`�D��=��|�z����R0�
D�H�	"$��X��X����dbr1�F��=�w4�w4WZ�
�����h�&G�ۙ�=׋ 脔F���t�u`��`����q����<?���åçq�|Sf���Kq��:ݫ`rƑzv싞ui��嵤�$L��� �o�@��^��[���}oۚ،��	4��`���*����Z�d�R]`KP�+��ը���׌%x���mz��D��2'�ɚO7ߖ��� s��#ВԔTBI[v�h���bs���L�=]n�*�������^0?��d͈��]J��Kk�[S��n�s�����z��C��n�m.�f�����[���e��͎����,�X�[�������C��Ǡ{��h��h���{k�;9�:�2L�1��3@�W�).�*����Z�.�.��)������^�W��ηs@��s@���j7���������k���`yIu�3�߳�ݿ��>�UR��m�+���     s�V՜�+�yW+k��u�y[ҷ	�	;n�e*^x�W��]��NM��+�6��F3�]���i��e��vބ mPw�{w���s��G�M�.⹺w��.�=h��lU�k�-�vs`�t�5�n[r���pM�f䶷1���.ܭ	e:�Y$�g&1�I�g�B�&��N���������|�{ܷ|��.�Z5�WD혘�h�7l�H��^��E�5��g�;-���4
`�N>ϯۚ����mz��E^�8<Y�&hu��=;��>n���,�(�'��&�bs�$AG&h���{k`}-x��W�{E)�Ӱ��vn��v�*����Z�d�R]`|�R�q̌NF8H�z�n�{����@��^��g�����p������:e�\��a�!����b�nY�7Q/z{<�k��Ir�n�m�~��m�^��^��~���a�ږ�.㴵H��X�u�
4DRP$�QS�� �Z�d��S��v�p.�E��
�n�>��`Y+���X�(��0l0HN-�ٟ�����~��=]���j�<�
*���Lx�r����`yIu�}�����6������~QUV|�l�y��&-�v#�P�M���G=��tl&.�7m0Wb�n��K9r��R]`_m������w4���	� Ln9#�/�ՠ}mx��W��������q�-�������?6�`u����up�t��D� BL`��5F�1��h�WAw}=�! ��L	q�0%čp%0.0Ć���(i�J$�@��"@�!)� D A7�1H�=4Ş��/2\0�I����3F�(���aHFe�8�8F
Ř2F�!�R`@� �`�q��Z��!3LZ(�܅bc0��vO�͞bp'1�J��.:SXq�4�B���5���`��f�{���'��)�+�s|M�P�U�S�'�|
����G* �]��qP�����h
��=��>נ{���^s�#����c�^0"���mL��_ZM��(�����uz�ڴ-����z�4�6܆�ey���+.��vT�]dԃ�J�8dRۅLx̒18� '��@��V����^0"��Z�5^�什\�%��[^0,��).�/�ՠy�U�!��djL�/u��"���mL��{	V�ط���H�\����X�j`}mx���H+ڭP"�TC��!��y��>�]��"8���$z�ڴͼX�x���XD%��T���[uv�g\��9�h۠�VN�ȯ-ݍ��e���;��Ƴg�z�ӆ��&?6���ŀ=׋ ���BK�mwN Ӭ�扎�����h��h�נ?Ss�y��9B�S#�bꚚ������"��`_u`���m�����.#=�&'d�b���j�=mx��W�������W�y.�!	o&��J��X�j�?~���y��I$�6Ĝ�'���p9   �  :����n�ti��i�-�04������v�͸��]�XS;�:��Ƌ��a��ܵ�y^��gFx�腎q����ۗ4�)���t7muu�`�Y��3]�wD�듪j�ݰ8pn�S��6PN��I��Px�iڻy�Ţ�]��vUvl�p�s3Ɛ�r�����pm�l:D3UV|�`������������8�b/C� ��f���DR �Rg�}oۚ.���j��w�}��{�_�[18D�Ƣ�4]��}����`Y+����ܐ�	��r-��Z��h��h�V��-K��"i9�qh۸��W�v����S�w&�Gf�9�nf�{��k�h�j�-�s@����HHI\8jt�u���a�\:ə4o(����wI��H�Q���j�/�ՠ[n�ء%�C��X)�Ū�����E����>�>��h� ��z�� �DB�	.��N�ذ�}� n���D�8�&
`��Z��h��ÒJg��� ������˛����%��J�nژ�j`[n��{�[[18�%�E&h�S�mLmx��W�e��t1m�V�Zz�뇉�X��̂z�9���u+q�T@���u��q������4|�}�?~�mx��W�v������w-I����@����]��j�/�ՠ{��:�1�r1Lm73@��M�>�>��ZB�H�bD!	��H��"āHD����0"ERH�c$a!�H����!H�`�!J���x�Z�����+C�䂐I����7M� �M� �x�:"y���Rg||Ll��	�"qh�j�-�s@��s@�ڴ}kO�����8Ԓ{lt9����4pk�#u�n�<��۝.ܢIQ��qh۹�^빠Z�Z�ڴ�U[QH�d&jn� �^,�
d���;k�p�Ŝ�)��S��SVW$ʩ��Xv�&�ژ��d��+pAb�"��Z�ڴm��/u��8AM,B��!�s>�ϵh����II����@�׌%x��mL�0=��ڹv�U�.��@���M�p>ub8ˌmm׮a�#�hэ��18a28�1�r21����W�v����S�^0%�e�n$�O���j�/�ՠ[n�{��q{)1�&�'��Š_m��m�J�nژ���e]]�EL�\�rP����� ��k�h�j�/�eUlQE#�I��`Y+��j`_m��m��w;~����` �Y���6Am  ;m� pf�˜�d�$lزV�);;��bV�=r�cãcN�Y�Qt���դ�*q��朜� ����W�n�//�sϬOv��`݋[K+,㭹+8�c{��wK������|���6�c��������� ��v��m�m]�غ�y`���7l�m�k�qM�E��$�M.u�^y���w�뻻��O����q����C\�Gm[�=��=�/u��f\�n�݌,�y^.{[�+��c%�E&h|��@��V�m��z�n�!I�29�}v��w4�w4]�@����4����;y0-���^0-�S�mX����KUaWt]SUk����wWt������ �Z'RPR�N	<s4]�@��V�m��jXp�'bJA2<�)���*��O7s��9g�a�c�m�L�U��}7[��sdm�l$n-��Z��h��h�V����+ ㌘LIŠ6�,BQ��2=׋ n��}v���UV�R0Y��4�^0-�S�mLmx��=��ٵr]\�*���`t(J{��p���w4�w4�����&LL��X�78%���~��Xt����~��o�_vyHנ�<����eg��`��j�N.�]��ɸuK���(z�sժ��wv,�Xt�����M�:�1��L�m73@��s@�ڴ�h۹�U��P&H'�Uk n�����6#�I�$�T		A�)�P�A6� �^,��d��ۀ�H�Z�ڴ��hu���O;��+D�]�utZ-Tȷ��^0,��͵0/�������r<a�[V�[Q�ӷn�7g�Ӻ*��ɋc�e.�C�^� <�\��f��a݌%x��mL�0,����:��cq
@K�L�/;V�}v���`Y+������.��Zgor`_m��e�J�fژ"Կ\�&���$#�@�n�{���>�>��K�*jHB$c"���K*�#0�*9	rB!#"`�		�:a$�c&h�f|�%���]�=<���,�8)���h��h��@��V�z�� �o4<N�ۃ�L���1���S�D�+<����],rƑzv�Nsk��,�L&H)�	���j�/�ՠ^�s@��s@���Ll�����Š?Ss�	(��9�b�9�ŀ=��:31"��L�A�0���@����d�m��}���U}�ݫ�Z�d�Wk�D�}�`�p�np:�
y�~X���S���fj�2�nn� ���zJ;s�|>�`o���I�TU��("���*���*��PEW�A_�U�EU�DQ�� �	B0T �P��P�P�T$	P�P�B!BP�AP�T �T"�EB#B �P���AP�� �B T )P��B"��T"�B"@T"0T"�T"�T T 00T 0��EB
�P��B
0T"��T "AP�P����T"AP�)P��B$B
P��AP�(@T ��T"�AP��P�BB�"AP��B�DT �B"@T �B+BP��B ���P�EB��*DT"��P��$EB+P�!P�EB P�0�DT P�B ��DT @T �@T �@T"�DT �����B�P�A` � ,B �EB
�B � EB�BB"�E���P�1DX�P��T"���#��PEW��PEW��A^��*�U�*����"������
�*��*����"���A_A_��PVI��o��y���V` ������^���@@h�@ 
  P     ��  P�n| I*�  T��R���
��H�U� $T)*���J  !R��J�@I �U �
�    ��@P)@ ��),Z k���R�����}ܽ}w�w*|�Q����o�Uͫ�����w�(|�����n�U�� ����w׸>�|> �z��l���/6S���jk�(Ӿ�l��^���cq�=�6�  7��@  � ' ��˾y�<�Z���[�P|�;�W��_^�<�U��O_�}�J��<�[�}����Wū� ���w�Ʈ��P+�^�sk�Ur�o]׈��v���W< w��N���y�z�Yr��V��Z� ||�@  %@L +�_r�B�/��� �h(YJ s��cJ�����(�[��Q�(� gE,�)i�   ���z唥����)K�p)J;�Ҋ�� s ��(� t�@�b �M RݹJR�ĈJ(
(( d�� @K��szݼ�Ooy�v��|�@Q�_Zs����y��v^M{{w����$�{l�]���}{�| �o'q3�vW�| ��Nv�g�������c��[}��{m;�.�l�v�}������������@�� *� 	��@t{��;���k�u|�W��<��z����
=��j�o��������[��m%|�$���]���� g���n��w�Y瀠{ԯy��חͫ���|��/�y��o�OoM�_Ozyq�nm�s�}��   ��AS�E)R@�"����m��E   <z�TOJM 4b'�T�	Q�OД�Ҥ�@h  DHCRTT` ����W�����/�O�k�Dᓎ��n]b\�Is����$PWJ���� ���� ���(�T�����C����c�F�x�i�4m��H��@��0&�$8�bF�4�
�c\���N�,sL����I
$����%q��80��4Cg/2�����H	XkL6p*F�1��8@�J�kL6p��)���F�3A6�W��o�����i���m����CO�HSY� �Ri����m�����:��M|�dj�A���@9\FbN�p�X9��	8�9�3�?���~����e��/���K������!-4I<3�3l<a�m4�)��
�h��|57�!�+�CF�n٭�E�RS.��ə�$|��{>�\����nn������#��l�H��v<���������y�>o��S���m�x��Ǿ����NX�) �(���BD 0#i��/<�f{�<˲z`B��npaL�5�N�����p1 pRa��a��s�B�&��a��n��9�I�]�%�ۜ(D��FM�l�rE�˭�7v���5�|�P��v�Æ�SG�sF���g)�YL���s���]ni��Y���a�����޷���$ ��o˿^�����~V�s.e�I�q��x:(# H5!���&�RX^s^s^��h��sɯ�Ms��9���~&$OU��
�&$1�m��2`���A��Q(��L�N&r�=B5I!	)I�i>�n�!Hj�r4�$)�.�HS5�+��H�f+��w��3��w7���+��-3�y�[4caҙ��[���淣���@cC3Nap�B����4��f��)��m�4xh�i���7� A�`X�1�Y�sẊ ��	(D�,$��	/��.�<ٳ����8�|+���׎�c��||`WF���R)v��*9�O��L|BB�x<k���g�[k3dѣf�Ѱ!sF��F�8Hk���x9�6�HD�WSц�HbM�]m$��_JSen��5�w37
�D�e�0)���04Ih�Yh�J��5�jFԃ�>��9��1{�Mss��p�[9�K�"P��7��p��tp��X���}I2#Ea ��_�O5�3�ǧ�D(b�+��h9�<�@F�!*K�eI� W&�a�(�,V1v���	"X�5�Wf��D* b:Cg
k�s�	f B�5s���G[�}�3S:j`A��R"T�}��h9�7.��4@�h�$T�#���q��a�И�k���y{�{[������cVXCi�z����<�A�����^J�kf�1�4��h�����h�đ�$��	p���#p�3�a��q�W4l�bq#sD�gq�%0����&!)�a���h�I\�Sz8T��Na�Ѷ��7
���c�`���M$�hф��hၥ��s���y�&��V`_M�`Ը��fuv;��~\�k?'����f��s�SH�)���K�_!E�^g����8fp��������������;XQ�S��O����4>{���1�8���Sy��o{uB�4l��rxB��kl�&�x��6I���F�5��:q"P0�ѳi�6h��^NB\��xh�8m!p٪�<��f�!�|��㤞�8rL2�|^C��w쎸A��D�4�O#.9�s�ik#�Mp�/���>���u��i��V�����6O�!	���G�X.��x�8<9���W$�pr32����'f�`zp����N[)#�ٞ�6B�{� \w?w��yi`Z�z*p�3�Ig���Ir��W�߸�hu���5$��l����B�	$�aYy���s��E�F'���Zd�RĠ{$Hƒ�s'8a�oY�8����S�~�׺��Ǎާ��j\�s�hަ�a�l�9�ޫy��rLi&!kX��0~D��w$p�!����P�k/d�icLcI# �-өw��&|�3[���hB�FHB��s���YR���ae-
M��(��0a�%��6BD�m�&F׌ڂ:���65�LS�_��܇�p`P�x�!�"@`��0Ӷrj^y7��y.y��ko��/ W�ė^�M)!���x]`���)��d!u�����B6�ÄB$Ck���ڄ����Y.}��o��u	�����og�OA�IB�I0�RI!Gp40(a���<����&���p4i�ә�r��4Lه+�fWd�p���S��@�5�0��W$#���4�0��l�xg=�G'�T�N E"��0J��4�S	t���˞��i�䷕�)�ؤ�a��<5�Я�|��A+�'�i��%L� �CĐ� GA�����T2BF�PSN�LӲP�r%f�C7�yJ_z1�� F���Y h ��p���!���i!VCF��#�:$�CN�;��	���h`ԆGF��&h�	���f�<%I��&�R.:�H�h��$bRi!��!Lf�ÁL(�kA�j����8$`�$�Ƈ�
i��X��3g$l�J\Y�p�0)4�ơ\f�#0ԉ����]D�Nk^y̷�D��׼�)<�l�!�ԄX���7NK99<���4�0��j���Sz�e��JaH)��.p�R&�Vtkt�8�
���i%��a#ɲ�����R����eI�ayL�'$ѳ5����֤�����$��i��L.�&��h_<v����,���6B����������NnRg"jD�x�0'�P�@3BFH&Ð�c�F��c$2�[s�D�����j�D�)�!�!��S�))�# r�@�d�k^�7�����q�ϰ%��!��/��nJ����k���h���>�C@��"��X)"Ab�1�T�5`Db��I�܏�(捜M��$Ja�a�B�p�k|���P�y颚<��`\5�B��f�@�4��^B�so�0ѳ��߼6zzH���H�&�iS4{.�=x��kf�I&�5�o|�ĉ�x��hy�~;5��<�Ar��zO� Þ�h���0ͳ���jm40�|B&���l l���L���5��.0m	h}�Ms�d$aS��ƛ@<�8B�����y�� Ad� �Q�"�$ �!�@d��i�8n�<}8$���6l�1�5��N���,ԥ�~R)�/��S��4;�fv~0�3���Ӿ2c���y�G$\��g�=ǚH]sYɽ��ӆ�ޏ3��7�l�!�7�0��F7�/���g��B��!w��2����t�yN�,-4o��q!4b�1p�ر#�9.:���� �z�.�c1�#$$l���4,d�@��d�20�4 #�@�6��@�$�ca��h���A�
�5�দ>�����Oy淣)�����8z��+�����^ɣ0ЄHA�P صbAX�ذ�"R DHB2��K$�D��	HB
E��E#2��!$	Eb$�Ba$ a$��K#0�X�	(@�kJȲ0�X���	F�#�E�	�jB��h�# ōma		�Gd��BKB�aK��0a�'��6��.B0ռ��!캺w�p�����e9���[	6V�$2MK�+�P�a���Jo٘�fK���94MI]��<7d�s<�$��9��m��֌����&*@+��)�/9�B��[�V��7O��$߇�^�P�$�����$f�=�I�l&���8l���d%0l����-0�`BR��s���Æ�0U#���BlDE��g,K����$��W�@G=Y0ۙg��=��ԛ��>_i��q��	�����֫aq���s�s��1)���a����0>��Ϲ�r|Vqo���-$r��-2���/m	i)Q�W�^ڪy�Ԫ�
ܕV�0n��q�m��
�U�!FM�e                                ��                    l�$�GP               m�Q�ݦ����9�<�Ö�j�U;<�gN�,@W j��j�����-�B� фU�cV�i�g�خN��R[�ZX6QmXI�6�i$���� ٫�Ά�	�`a��5�<��9b�Z��OieZ�VI�4� ��xm3[u���i����I& ��|}9\c��9�vWUpR�ҭS@ �[.��k.���L�ok�aq30j�`�
ۀ       @              H   [@ [@             $               �                                  :���6��FoY,�{Zٴ�R��� �n�"�M��m�6Ͱf�v� � �i���&�JÝ���W�6��NQ1Ͷ
0^���nϙ����4,p���HҨUhʴ�+B̛��:C�;m0ݲ�f�ݛl[Ce�.`� 6ͫ`\�:P$�k.��ͩ@ ��� ��:�$���[d�g?��o��\��#M�[�2ڒ�< A��5,v�*��͛� �Ym�]"�6׭� 2- z���H1r�;fp+T�k;=t�֢ ���tM\;e�$6�߯���<!�z������9��im�.� k�;��Q�V��N�Y7��qR҈m ���R��ˬs6p���Șh��\�Wc��UBll��c���yv�eGJ�U])-K̻�ӰlIm�yV�Ԃ@ m ۤض���e���9Â���ֹ6v^�rP �;jY$��ڭ��*�p��3]<����Ż�m.� kbnPm�/p��#��L�+�q��Ut@ �Tx� [C��5�Io�\��[QF��>o �R�]�lc���a�]R�tP][]�j��$ �ࣙ����% � $K:�%�n,�*V����j�����H�Vhp[Knݥ�m�H�"M��r�ܻ*�6��=�����j�\�S�m�e�8�[�᪱�[G ݨ�m��hm���%��`�@�U�(Mr��6�PUʯT�f�ջ0�p� `(����YW.ݶ�[N  6�   �     �$    /Z ���A%�򴍶�U�_=�9檫�����V h:I�F�ݣ���� m[A�lh  �l��t��a��`�e����ږ��|�\��'G�8:Z���ʪW9~���'`;v�.�zh�3�m�@��gg�%�l�R�ў�N��w���Vy�Ú[aC�Ύi�y���9[���s�*���=�,f"���c�[s疫�C����

Ut�T�B�F���H� m$$8�mF�Kom�Ŵ&�g�鍶p l��d�ڭ��N�[\[x�{^�$mu�¦ی��� 4W 6̥I��,������h
�Oh[iP݆��}����d��ņ	Ҡ�V�������������q< Jp-U[)��oi�A�[{5�� :U��]��U�������I����)�6Z:�z�H rI:Nm۰���`�s��`F�kTq��}�  UPU@*˱�:֫�ݒ�ڥny�M��Z��mֶ�  Z�M�V��3� ��tJ�� ���Ijc�ݭk%�i�M6�� �(�n&�5���r�P  p�M%�t/dI��Gdx�+I��²�*��ͺI9�ih�h�[V,�L�����x�-[%��=�e��)G:�ͪ	��	"d4�ˌuJ�M����:�` ���� �U��Im���*�nʮ�*��R��WUZš����   h�H��m��l	m���m�    ���  h 6���&�$�հ�ٶ	.�¢�)_h�lR�jt�iU
孜��#qě-mU\fבhe�0v��@�Nͱ��L��m��  
I@[@�P#]�   	�-  �խ��b�-�������,te�Hsitֆݱz�ZRCk%��6�\Ɯ��Q��z�#S��U �m�2H��t�.J��5Zm��m[  m�ٶ�9�MM����y��rA#Y�Nn�@ �oN�uOnܖ�p5�A*U���pl-@YF����:��,�S����U�WHn�@AG+*��h m����i�b�U[\��Ul�J�+��dV���
��ļ�+�9�hmu�-�5�[%-����0��zFFp�%�P媠 ��\vi�4P�c�܁�����c�8�"[v�`�&�M��f����"� pE�����%�3�V��4�m��$��-!-l�i��=��#���kD�.Ꝙ���:T�Z��&WjuOJ��ֺ��� �!<u��oP  W-�[��m��  �q6�a��^���d R��m�m�ڪ��L���]!�K��l m�l�   ��� ��6���~�� [@K(�@{I�� -�( l -�8�&�fۍ�d� ��mn �Im�nm l���T  (8�"�;EǕj�,��Q�=*�T�I�ā�޲Z�L/O�D�6��1mu�1l��
 ��l���$���I ��%�y|MX6)�!e�)`:���j����a���
�8�Nsɩ���4�5@mN� c%U�U�N8���+j��BsgZR�  t�n�5��Y&X5mk�C��Re�[#Ci�j�%f� �`  �m��nqm�K�k@�`/Z9�ڝ��^�E6�D   � O����  �` � �  ���6��6�&�]7f�I�� ml��m��d�-�M�t�;Z��[�� 	 �$  � [@   �        �          m� [E� ۵o\�4�2m�� ���L ���  ��>��{k$�� [N,6�H    ��R���|������UTZ 8�  �6r@~�O�����l�����N�Z����W`*���(t$�PM�C�-HFf�n���VV�h��3�u]K�&���Iu�%c���	66�@[ �v�p� �	�__�_�� m���  8�z�F�ݲ�ån�� �UD�[@m [@��-R�UJ��*��K�z��@i5i0�Y��W;��+����Շ��� n�����m'`6��-8-�m�6��%E��az6�m��N�Z�W�[,�3��X�֖�e ekj��P'�E[P�m�[]#m�A�@�m��3m �d�$
��M�,�U��ev���M؝8���`��X$I�y�*�K��@U[m]!e��56U5.mV�늃�&Ե*:H�c��P�q��mml�[�@ۘ���=�9h�A�`�)m���˵@[u������.�hK݉B�t@5UR�]�^vn�W��V�umHm�\Ԡ3��5��矾�Y�ںڠ;5J���j�ڐrf9t�b1���j�q�랠u/#�d	tU*���2�S�'m�֩��UP�V
�5��m�[n:��%b҂�Uɗ^k�y�tl��-��<[������;���*��PS�ZI�6� 3��.�%p;V�u�mPq�A�C��m��`   ݶ -�m� ���E�յ@+*�t mUUw@U^��L��uu��m&�s��ݻbF�(j�� m��@ݗ�]6]�^�e�H [M�`3���J.���WU¶�:�v��vٝu��md�m$m������ֶ՛a���t���5� 	��K���lI#A�@+�ꭶ�U*e�*�UvUhZ�iBݳJ`�تt)2KN�ЋP�8X�1t���U�#;��	8��i���ܐr���K�N�k��M����j�n+��F�@Mk.�  9�h6ͳm����z�l$	�HV�6� o8��m�a�\���x �e�%kl��r@	-�G�bK���.�UP!��uu�ɴY���[�nHEM�!��޻K*�H-��	YYL7��L�B��J�	�UyeW@�D��mK�
e{j؋*��S��l��+�]UR�@�UĈ��}��X��f[! H��)nP�t�u�jj���  p        [@          ���                   ���5�����l���@x�x���}��V����9_u   8���ֵn��4AU?ʢ��DH'���E��!bDXl@\W� !�&���'
	��P�1���|*�&�>V�4	�O]�x�m��h+PWjb#4 hT���F$H1�D�ŋB B� ��ۥ}�G�B��"�]�1�$bĈ�Z/����"0�	�<�D#1�=S�p�==��`�� E��H"D ��
DG�T4��
�b�,8"CbW�h��Qҋ@��1b�X��H�@��!�x�1a���"8�~> ��؀�-�F(�M�"E�>A_ C��` p�"��Aீ�E2"F �"$b `
�H�Sj lAG@!�x �]!�� ��t*z��j��@(A\PS�>��H8$X	�0��$N"�D@�0q�J�pDH������>C�0}�:,�z"J�4����`�Z($ت���t@�)�*�@Ck���E�}X,��1P�hDb,S�� >�@ț`DU8��E U|Q�">��0�� !@�`�&a>,4\�!=m��#[��     6�   �ie   ׶�=;SNh���pl7n��ڂw]��mÍ�`�	v�5�ڶM��Y,� [@  �[@  6�  �      m���˭�f��h�Vvٶ�Z�˳��l�ۨ�\N��m�"M,�w\��V��Ӹf�v���#̥�.y��Q&�x�+�4qWGm��'�����f�&%4����bkgh���v�^1�;�
W��%+f�/@H�����C;�sT��q�E��>^N�ٓ$ E	���l�'�� Njwh:#m���=�j���w+c�9fC.����o:��f�mk
��$�5�!5Ι�ť�Q��,'m���*)#�ܡь�Jl�z�#�:mK��Zh��&d���Z��˥{6��V�)�l��ȁ�����`�	�!Hj�݄��GK=���v�]�hԫɪP"�����k:ݝ�]I�)�®Z-��b������gY�qe��j������YE�C�.6�+�p��l�	Ә1"i6x��U��F���hV�\m��Ԭ��;��:@�a^V�8��Lu[�{v����T�H�h���}][f}j�!��v7lg��M���r-*�U+�m]�<��9��G q=8m��   $�"Ӥ��h5r�67T�)���c��[��͍،lpOYT�K#uY��������k�g6�.�V6��8�kW��Ƥ�K^�v׎�nt������-�6�'��,g��ҦN��y�N3��W��s\e�+c���8�B[�N��g��&�6���e��Ƹj����4!73J�pq��ڎ:ԗW[n��+����W���X*���cF��A$�+��M;)5�iы)Xݦ��y��	����"��s�n�T���^WR'F˺&mH�im�`h    ��8��G4Q_���>��{�|@�خ*��4�tS��' CW� E�(�*��A4�(qG�o>�#5T�]�K�J箠���m�� %�#N�K{+�1X��t���7[%byp��CM<���{n)��vu�ɝ���ym#����	�!�UZ�5�m/�V�[��Fn��uw�u�PO�f�us�C�@M��n�vq��%0�m7<���I9=;��Y��ӯ�A婶�wjѸѰ��swR��7W�#�mG\�).e�$�2\�$��%���ce^p�3����vpbr�2F��H4��ow�ܴ^�� �[2��n��-���OV�@*�W\�}l���X��Si!	Uv�^����/�� �l���@�tX٭��xkO5�/�� �l�]��*��=�T��4��a����� �U �Ҹ�� g��wM{�:Y��(��]Zj{e.U��-M��E�C�n�6L�F�\^lm7}���ZW ��d�� pr5"��� �x��fUĳ�O�������F]�d��2y�P��Z�ڥ�֋K0��� ������\Iq�l�<��=0��n ����@/[2y�P
�+�_[2�뺄��d�I]� ����5�W ����� {�կ�h�g
ڷC\=#h��WpWl�Md�9S)+sBѐ�,r�D�al����N;m��5�Ҹ�f@=m� ��P��,l��%�m���� ��d��@9ZW ��Rj`4��hXj׹y��lܓ�߮�'>W�v(���p�Y��.	MՍ�7��a�rq.(�Ǔ`8�2l��Xw�@��X�:��Y��Q�,�:���w���Y�
�W �λ�س�Ow9]��4�/�z�tܮkS���Ӻٺή�_7/4q�U(Y]�����E���o�@=z̀Uz�+�p�[�I�0Z���@=z̀Uz�+�p��,��u	�!��*��V�<���?lė%3��Ձ�Z���-�P���m��{�f��ŒO>�훓�b�b��UUs���x��v�H;,mDY!foY�^� ����+�\멵?]�MT�S������{�nM�WH�5'\4U�`�ю;`.{�l%�䬘�/�{Z��8�=iΤ�@f<�`{�y�F5y(��X���&�}�\޳ �f@*�ȸ��b��1=P^�\޳ �f@-}^ t;��%���Z%V`��X�Y�_U ���/�n�!�K	�V�{��.%�z��k��ŀ}ė8���/���e� �p�l��ƈ2�m �`����e5�r�Uۣ�Q��v1�v�h8�]�v��J{pR�������k]CEcr��8��p�5Yi�V]�h��u�1�sɺp��3Ŏ���M3�utKEu�������Y��oSh�V�K����ݳ�rv}�����\P�wNzy�����AE	eB��Ly%�F(�BگS*��\6�w���������G6��rk�	���B4�׵��M;q�6�Ȗ�^��yɮ̍{	]��ظ�s3w�o���� ���-�2��d ����B*^8�������%�6{��X}�ŀn������F�u2"��\޳ �f@-}T��W ���5?kthXn�� ��2y�P^�\���d���o��n����r��f@=z��7gd��P8;k*��)]}9;6gY'qsݗ�L��\ٵ�wHfX����V��)ȷ��OT��W ��d׬���x���p���R�J��7{���EC�%D��Af�J"��?g��o� �T��W �e�Ě�oXa���׬���B�J��ـo��Xۮ���IT�ʰϪ�r����� ��2 }KM�B*^8������\罾�>�������vz�����ѯ��y4��kaw.��S����+4�1\��f�6�T�[j	i"���dE�+0��,׬����r����Z'�z�+����qg��}�?o��^�z̀_qpIM1�f�z,�@-�߳rOo�f�ERt�{��6���ŀk����5yHܳ ���/�� ��2y�P��['	]��+D��w�� ���X�����������mm��	#�o=�q�E��l\��Þss1t�GBrL8n�ف�����q�K	�W�}�����x_ul��=��,���vu2J�������r��-�2�l�����&�c��;m� ��Y�[f@-}T ����KZ�D��%T�b�ǟ���̵`7>qa|P���"(H"z
�1w�2���]�ǜ!,,�� ������ˮW �����v�qh�����:V��!Z���۫[���mg�ӵp��ڠ�����i��m�������p�f@=m� ��*�VF�w�M����ٟˍ���,���`��xZ?i��%v;aDJ��u�2�l�W�@9u���n�7;@B�Ձ�s��P����7�|���ٟ6����������!��*��W�6�v�3m�n�>����q<m��w~_|�{�u@r�m��<)��l]OE֛�� ��N�K��W�����ˇj�z����X�6컴Ӥ*N�x�����.��m��U��n�Cm��l���P�24�ղ㛜O(�sNl��:t���z��V�1E֟�>���'�m칗��Pf��
�N�ΰ��97�=$��>���❣7`ܛ�O�:e{Z�̺љ�b)���9�˗-��ѹ5e)�k%����9�z��/d�z���ֲS0�v֔�]�/lW�5F�/������Iuvb�$�m�>�$�툉6���$Q�L��BϾm���O?"�e�����[o��wf���}>�sK��˨���X,5k�Q$��߳�o�w����I��=>����؞6���5��$��YW�6���=�1��������Iuvb�$�z��|�UЪ#dj7yDܬ��}��g�6ߒ��_|�Ͷ�����o�w�����Sk�v�p��^<]w8[E�t=g��=Z!뫚C:�Vg��̡�,m�VvI��nէ����?��D�^�~ϾI.�b/����{�|�\�`�hEr�B����������� v"A$ �` �Cv/��$��?�I.��Q$�֩@vu2J��U�ͷݻ����7�ϾI.�b"I/^�g�$�����x�D�	=��Q$�;�|�]v�D�^�~Ͼm���Om��5H�v:�d�|�]v�D�^�~ϾI.��Q$�;�Ͼm����Љ���U�ە�T�۩X��Ű�ּuo):��y,�)$����Xt����a�޳�_^�g�$�Wf(�K�⿾I.�b"I+�.	7��f�Z4;W�6�vn'�ܒ7��z}�mﯱ��o��~_}��qI������n�S��{=���6�v�3���BKQ�p��R�sZq�CU(Z�J�`kZHͲ���6�+
F��a�*M�,�L��8;��Bi�F�H%V#Bh�b�9���Y�(c�m�� F��p�ќ�2養i]��v�at�1I�*BCY��y�����5��49�N�A��o� d)D�z ����� )3!G�	�zu�!as_E��(��9�$��D�$���
 ���@j��+�
,Q �Cb�!���*i�x#�`AO�8��� �9�{�����vb�$�R���{��7Rr�}�o��S}����o��|���)&�{�߹�I�t���q)#�z��+)-f6���/��RG������i��/ߣo}}���}����n+UdeV��9�s�^v���&�af6�p�bې���+��D��U=�̸�~m���'����u���b"V\��L��e�oW�����dMQ�x7-�<m��m���|ݿw]ݛ��������-���v]�G��Z�� ���E��ȋ$,�������c~���w�9xf}��˻z������[of��d�T�"+��=�$o��|���~�weݽ3>�zw9�n�M�!��B���@�C��"����=C���w�7�\̷߿N��>�Q����_|�{��O<�$������ͷ���c~��{��l]��Һ�8��$�p=j�=E\c=�Iz#�N��;K��#��P��d��Jr���}���b�O��+.��3>ǟ��]��Fl����H��{����ʥh�Y�ͷ���c~䓾�|�����؞���VϾ��>�n�@AaP�%��o�~�������_c1�ߖ��z~��{��Om�����d�Kl��o�w����r��I.��Q$��_��=�Y���7\MQ�x7-���og|�>��G���_��m�~������ݛ����ED��%� cD�D ��{���_{��ߟ��q���lFt�B:ڦ�d9�  K6��µ�x��YЖn�]<i�WH�y.I�#M1�� v+Y�ܶ]�Ѭ�����#�n���Q!w�}�����]�\�-oz཯J9MvB�.�m�Y���&sc���lB��Z6.сݓ6]ےᇛabz2���gos>���&�N-��3:M��8ȘF��{��^�Z���w~��Ē����>��
9A�\�m�i�����r-����퐚�I�@rJ�]���7c��8��ͷ�鸞6���ߗ�$�]���IW�+����&F`�����կqD�^�~ϾI.�b"I.~�_�$�Wf(�J���m��cY�����|�]v�D�\�r��I.��Q$��_��J�D`kk[�LI�"I.~�_�$�Wf(�Kׯ���%�lDI$��h�v�U�;U�|���q�۷� >���y�����ܶ�sϏ�|�޼�]���9e��p��G
ږ�@��;=L��(�gg����d��r�N@����\��"ҡ	�T��o�{�/�m���f6������$�[1Ē_Z�1-��{�Z9�m��}�7򝝰��TR� T!�Q*@V���-�wù�[o׿l��e���t˖��Ț��x7m�<m��|�>���6�D�^���|�]]��I%nU^�x�ַ�b֞k���ldI%�o���%�n'���n���ͷ�wIA�[�޲$���������Is�ϒo�w!�m��n9��:ݱ�(ՑÆ.nr����T]��W�3ڛWd�+��4��&����E�}�m�n�1��gul���l������䒪�Q����r����;�g�y.$�����d1��}�|�����q<m����)l��+E�Ͼm��܆6����/�s������1~��̒urb�$�����$�����N���]�����ͷ���cm�����Ϳq)���Lm���y��D��U-v����n�1��guk���l�Iz��@<��Z�-�F�$���C�+��f��t�Ib15����ä5M�P�9x�il�����mX_ul�9^��l�^� 늭��o��kO5�9^��l�^� �M�ϺH�	�*�2"�,�?n�d�Y�V��9^�}�m��o嚱k܀u�2����p>^�4�T�L�|7$�t���4����܀r�k�r�\��Xw�� ��d��P8:���Ӫ���Lp�^e�0n��N��]i.�_1��9v[�j�A�-uJ�� ����;����f@9\��9qn�<7M����ͻW�����VGVd����.s�����u��*d�K]� �nZ�=76bID8Ǔ`<̵`~��[�
�x7m�`z�f׽ـwwq`{�$��� {|���(ݎ�A�x��9^��ِ�f@9\���9H��-�����m��j.�6th&�Ͷ�$
�U ќ��;��x�4��xy#��3R.���Wz鮬Kp-��&��a�l����N9��yyGW7m\�<�<��*e�R�NjNފ�u�N�wϮ#.z�T��HR>��l݁Nޥj��\J�4����Q�5���,x����t�z�!�6�vct�It�80㞫Ywfѻm`��Q�e|�շkZW�!�
�
j��f^V�Z�����������:9�-2�Df�|����%rm�v���U�U���f����ŀy�ڰ=y�ܥ�A�<��&f�f�Y���^� �upW��u�2}B��m1�LI�@9\�6��͘��x�Հ�� �y�E 햺�h�ـu�v`��,�� �up^-׉?��-�p�f@:�2��W �mpy�G���a���6wg�kGJp]Z�����*��b��b�u5ّ�cOm���;�� m� �s��r��^� ~�VZ܀VK��e� ��ݘ.~❠� (B�2�E"P� 	�WF���}߻� �����ײ� �䃲)f�ḿ��j��\�"fZ�by6}$[���ȋd� ��q`��X+�\���/�@�s����f�Kw m� �s��r��zِ��K��vÊ�slIDGNNIgui�vnzu�.�#t:CRÌ���Hݴ�z17� ���9[\�l�[f@��6�A�#���� ��ٞ���2Հ�2Ձ�k�lGF�TA(iP�� ���Xwwq$�K������fI�磀r�\��i�x�o����׹b�o� ������޶d�R��I�5	n�܀y\�6qqq�fO��-Xmڰ:��L�W��&�Givk��=�����]�^--J�-]6�"��u�2�tM�%�ļ��9[\�l�[f@<�upt4�j���k"-����q`��P+�\���/�@�s����f��@:�2�s������zِ�DkH��bor�x����nI�}�r|��J�d�(Eϯ���R9V�9K0�ݘ�l�[f@<�����{��������{6�r��+�7/l�+QjzB�x�����V�N���ZT!;l�?~� �l���\���>�m4o�ſ�{��n��� +�pV� ��̀}�\��6���-׻���+k�{�f@:�2 z��m�ַ�b�ٮ���� m����'�{Ǧ݇���ZUl�6}�j�ĒO3?/�v3��ۛ�aHִ�1��
եeR	YRVVV$e	B4|C�y���k|\���0d1�B		4`@�@cN>$k�dJU�Q4@�#˱�@i���W���2�7�@��Mf�6bbI|�&��޷�����	��#�VR�I�JJWMS�',�8��5�H4H�(����E��"x�]:i��� rp�3iby� /���HOR��(F�*B�(J�X�jD�
��+
¬hB�
1��F�ynChB� ���X�>;.m&x+�pT8@� D.����If̰�	����C0����2憙��Wg� og����-+�jP�(` ��!��>LM�#u16�k70���       m�5�  ��onִ�0��5t���V����rN�m8�ʠr�'ok�C\]��mۀ�  ��l     h      3m7��-�w]1k�i�c���m"^�#��/=��������6Kbٍ�Ϟ�����@��D�*��um�'�"n]��q}�[��8䱟 �[���8���\�[F�/���75k9�l�N�笨�ݘ��r�����2�=���NZS"�j��۶�0�`m�B@ 6���-�Ś�rlpNP
���t�a����矾��9��m���s�P�6��ە�n�WF�,����:����B�Kpb�n�nJ���j'��p�3#�F����ù�'5JYn�=���x���"�
���{lKr��z�9�$�T|��O��f�ٕS��#��U@U]("�ftK���;5luY���A¬j@�Ȱ �b��p��W��᮪��{XBy�x��흝�zK�%���k!ur�nY�Ō��٨��9�kv����o[mà���6γ�Ij���mR9�%�zAsذ�e+ ��v,l�6フSm
pOh�T-�(��lh�mZ}v)�c����E9�۫m�;Uj�a��+U�Űd�V����	�YZ�%g:�T[5^86Z   	5h73��:հp5HKhs�Ty�nzQk�[���(�Gc�j:Ӟ֩� ���Jd�����t�΁�W���r��k]���������m<���-n���v:8ے�s�0\uV�ķV[t؊8˓��v��Y�탊��I�Ǧ�VU�1v#Ī;�#u�M�y��&��+���:��[W8z<�����]����6��Wf�OZV�A�K�Ͳ���gU]œ��pާc�K���9����1��gf�q�
ݻKi����7)�����Ӥl��s��Um�Z�   N������C����
��t+�.@���*"|��X ��Gj �Q9�{�k� ��1�jӚb�m��Z� Y+�{(yZ]�ض��ٶ��q�����\����|||�8
���l��TX�/F�Sm����&|R�xZ��iݬ��C�r�k���;.ypg]n3vŬ�秨oEgv�^ �URe�"�5N��v��v��a0�q�����1�tu��#<�|����Lr�{{:w:�FUV����w{�׻����u|�z���]]�;Z���N&�t�,n�~?w��f�'O]^�q�E%;`[�g^;Vj{�m�� �ZW �mpwY��D`kH��bor����� m� >R�m��QȚ*lCnl��՟�fZ�;�� ��n���J���`y>���fZ�?Cc��9�6s"��g�;�%V�Հwwq`_��z|�{� ���X_��7"����-���C����\�7�{&�&����@�n�ҙo�������[qd��Z������^���l�[f@�-k6-o&�rOo�}��i.
��c2 ���<_�?sٮ�7$�疬�c��\��Jdy&�&�"f���(����nڰ<۵f$�=�M�����7���9ƫVJ�=Ğ�3�=�M��m͆%y�����ȴ`kKQ�bor�i\���=�̀u�d ��;�M[��F���e���s�&9�0&�;V:�� ��\[WE�9o߽�ŦQDIv�㔳�5�ޘ����<۵���Ky�vA��`d3v�D���'m�����$�f��ŀu�Ǧ׻� �u�)'#/#�Z[V��ٹ'��ٹ���TH����T�Pڢ�C�?����f䟾��b�>�����^�-X�s����._�M����M��7jëV�%Y��@��A�l�7c��vHY�~}�{�s�3��<ݵ`v�Τ�
e��B���a�VW��2k�V���]���·�OD�ª5,�Һ�-���wq`mڰ;�~K��9����l�~"f�(��
�T�+ͻW���G�́���`w�ڽZ�ɯCb�ARD��D�+ƭٰ=����Ȇ�-X=�X�?i7�GV�8��K����m���`n���ͻV�K�.!%ÃH(��#��S�M"x� ����s�ܓ������p���HB���ͻV�qj�����g ��ـw�w+R�T��2�I[�Sk�t��y�^!�V�v[�&wm��s�]��4Ԝ��I*������ ��n��[��\Ի!��j���U�A��&�DUMR�=77���2dn�����7���s��@����d�,uB7dR�#wf���`y�j��5�6cɐ�&f�QJQU3Sa�����J�>���߾�Հu�:�ռ\9�9[�6�h7�D��U��`y�j����Y��27vlu�Vˉr������S+�_���������6&ɭ6u��  $�$l��fI�Ռˤ�s�,:����k�tv�2��7;�u���;u�v�C��ͷ��%��N�3��M֡�YN���;l�b:wO���>����H�B����}9��t��4�Z���Q�&�]���f��b��P�G�tVֶ�s�ӹ�eyzۃv���e��ׂ����s���U�����B��bWX��G�P^�lE�ԾulqF�W\�����V�설ab	AQ9*��mX����v���������֬�����Ɖ#��ZdV��wf{��c�e��e� �^u`zn�H�@��HB����nՁ�ݫ>�9ū�dz��p?���}�]��9��Ul����<���؞U��m͆q(~�����喱���x7,�`�]ۀkݮ޶d�f@/�X�+� A�v�9��Z��C�ڝt��Tn�X��7�T4T 9)%�H�e�A�:�v)o�y�ޛ�nՀ�v�~�=��X�XB��I*��"�,�;�wo;Ép8����q(�9�\\�\�)��Vּ��p۝�Q�����[��	�M5Iu�rM��Vּ����rgcwf�ǻj���TF��n�or z�]�Tۛ�nՆ���wwz��-���D�*�PJ���nl�5%�w��n�ڰ��Vz��5U5H"�UXt-��<��F��Q<�����Z1qn��n�9iT�@�jhVZ���ŀn���ڻ���>a��z`��}'"��M*���`6ݫ��j\��6��ݛ��q`~�VZ�W�nYj��ë�nl�qB�󉤖.rm��V��ŀ����n�T#n�[������v�vl�mX�j�x��=�ˀu�xj?(IT�Q�f��w��ff~_�;�ʰ6�����%�$�%lt����MWbZ#5�v,,������7!���� �籯�_��̵`��V������b	PQ�U�~շ?�I$��67vl�mX�j�jK�!�1ljP�b&)H��UV��́��ڰ�d ��.�*�n����a���Ż�a�I(��~Vfe� �֝X.O5!D���D� FH�@�!��$D��V��B�b���C������������I�R�IU�ڰ��X��W`[\��2��˯�h��K�,�s:%�Y�zS�)nn*��CA�V�ų._%ĉYJ�mW�nYj��|�V������\\_�33-XydFU���H7\V��vg�l��`��� >���:��5�$�ҩET�M���Հ�v��Ē�:�eX~����ۙȆ^5Z�U����������U��6���y�������(�
2ʰ��ۀk�s`w�v�۵`Wq.r���"8$ Z!U�`��V?*�@?�����s �At٦�\�*�m�� %�/N�h�3t�cN�]�����s�����9��T��A<yT*���U��2���cm���(�U�j즞]���tva!�>���\v#\t�a�=���9��Z5X��c�ɶ/�F����wf6�G��y�n�{m�X/Pmc)���Kt3�4l"]nn�V�f��w���Ը��IR�5^9�/JOl��:�ݛ���ݧZK�S��[�%_�q.\x�R7PTU*�cٳ`w�v�۵`�ӫZ��u8�p���� ���,�s���K�d�ݵ`�[V���q.Dy�E9�U)-X��b���n���� z�&�������'�w,7�\[�$�}�mX�6}�j�W9�ũ$�ww��5��ک� ����S&��k�{�̀[l������$x��e��Ul��)`8��)���Y�nFti��jlM� ��\I<��y�,*��UL�����۵`lu`5mp{��I��o嚳[܀[lɜ�IZ&`G �H� �	H���&	�%	p"�b�%��B�Y���U=D�#�R(;�z��̛�n��A���/�a �
2J����k�ه�%ě��ذ{�ŀ����MH�uARh����s�v�vl���۵a��M��=p5��u8�r�TBvـw�ڰ>�9������6���=���s[Y��y����ݱM��b�Նvw=u�(V�6f-u��fF����-ͪ�`6ݫ �MՀ�:�9��f���,�R6���,�`�[�?��ų&��́��j�m�V ��C���,uB6�R�^����Ņ_�8��"F#���@���Z��	��Z;�*��L���(J�@�qp�����,sB0�p��g�ˆo����D�S�zC��a��J=�'U��� ���{��S·���`A�eBP%c��)5ߒY~�\e"BP"�16p�\Gĥ^����$�ٰh�,��!	 �O��
�`e���(�*J¡
$>����#A��,���S��8�E�_ \3��]�Hh%+i++$�`Ҍ��<�۲!� ��{<��� x�~�E:�6ն�Fö� ��BI �b� �/� EA��.m
�`�"x h;�X & ���#DG�P4"�(�A� �����ٹ$�����Ѩ�
Ka��.$�}��V֛��\QܬȰ������7��X��@;�̀r݀}]��ِ�[A=�LZn�q�Q��٩�k���|s�;�.�.6��������w�ffp,$AFIW���\����n֮..j���\�=A��Z�_��I���P"��l�xww�yڰ4�^.s�Ӌ��6��R�T
�*� "j,��V��j�<םXl�xߵݎ�J�%R�*��Is��qs����`�6��[����$$V,# �|�@N*s}��7$��YJ�mW�nYj������[�$��s�\���ﾏ�o֬w�Ձ�K�����r!9>En��+�#R�՞�u�룑�����j�s\$P�meL��������X9Ö�Z�2�eѓ-��5�d���?ʀu�2��2��W �r��),-�C�׀w��,�9��s���8�.L��mX5f́�ϜX�1�E"�
�T�w�Ձ�k�l��-\�I|�%��O�ߢ����V��5���� ���>���w��a�\Zqs���Ǜ�`1l�P�bf+�7\���zِ�Y�+����Q��bՂ)M�� �����v`�|p�֤�t\�t*Ү�*�Tb��c��-���ܙ�uӸC����v&;aq���U�4YM���z�n�ʥ6���j�f1]+�Y[�eK����f��Gm*g��Nt�&����'I1�����V0u��������cgsn8�&W�]َ�ƞ�rvƔ'v.��6���]��=��<ڹ3�u�F�޺����V�]�{��w����ߜ�G5��T�Wgv͸ܣv��.��gcu�T��!�*Y��a��ww}ݻ��ߑq<�TEU 5�ϭX�ל�l������R�IT�ʰ��x��Ԑ���pٰ=��zݫ�C��֧���M���t�r�T����l�|���[�`{�v��u��E���$,��\_���{���ڰ=�;Va�s`zd)�"��*��EUTX�v���5�foW@q�l���˜�7�$O蚪REͫ�Z����Ed��Ok'�����^�8�͹��Xv�Y[��4T^5Z�����`��s`~r�|���qvA��Vn��|��(�*�?=�*����8�s�N� �
�T>E��<���`7�Ձ��ڼK�Թ�*�W��!L��R��M6�w�;��Y�\J#{�ŀu��� ֻݮ�9y[��X����Ė��#�^��T��j��^t��׀}��vH�"�H�N�j�;�;Vˉq-\��8�>_O�N�{� ���+�ȥ#*�Ke���\	���/d�l�E;��EX$V�:S-F��ge\w��� >��n����?~���8��#��<�V�dF�L���jH��O7`W�@=� � ޹vf%��8�<�����RX[�m� ���ٹ'�{����!�Ӻ@7'v�\}ۦ��Mr38�Qx�Ӳ�I|�G8����=[V��e��u� �B�fōn�S܀z��$q/n~Ӡ7�j��|�X����Z+dM/,��%��1O=�P������A��K��V
��9n�R�@U*���2��|�X����d=[V��ҩ��DUP3E���ڰ=�;V��:�??S/9ż8#�)����"��U#�v;V���d ��.�>���{�f@/�ri�څQ1\����V�s�h�93�j���lܓ�=�f�(�A HX�0)芔��)r�����om�F�/#�+p��L�q.!$�����mX����I*˓c���uB���a�>8]sڷ�.�κ����ɞ��KH�ѧl��t�O����2��\ ��]����ϐ{��� ���F���ti�V���0�ڶ����}�j��Z����3t6H��AG,� ;���p��L���,��v`�ճRjG#��U����Ir}��K��V��s`�ӫZ�t�PU�h �x���X�ӜIe<������8�)s�{�??��=�� <�͊d�r��Z� e���v�EĔmuW-;#�d����x�&�L�]g1:��yܳ��=k��1�J�ݡ��Of	mLu��`iZUAA%=7��uڰ�"�2Y���:q�χ���\0`l�i��J_��-�n�5��=l�'��.5��ݪ�؅ɫILrt�@��GF�tj㍏&�r�WR�\����Y�����c\��ǎ����t�-���#g�ll�ne�^|=vJ����l�Zu`~s��$���\�y��zj�*I!TLW""H�� �֝X��Ł޷j��w�o8���s��S��=?�j7Iy�q[�w�{���[2��\ ��]�r�LMVcz�ܘK�kWr�E�0�Iw�}�`lf�6޴���$��O"����#3���7j�:�wf��K�s��B�8�-����͛�nՀםD��,�%wD3�WP]�Ƶ�@�9�Q��s;���h�0�sdڜ{Hd�k̀w�:�?C��n�.s���H���d2l��gR�31J
�k[�r��ٺȑ�N!� z�7������d�/up/\�VwihEAV��0߷q`��������)�v�����>�߿�p>E"�n��eX_���??�9�?C��9ŨIqs��7��צ����:�pv��zl�>{ݘ�Y�^���X�*� �=���
G+��rX��^��h��lk�6H��.�fF��)� \$�r�2�LӖ[�ɭy$�nl��v�G|���?l?
����D9m�����%�q#���d�y�`dn6�~s`w�L�|�R/� ��ݘ^����ϸp@,A�HB�%`RRPk� @���B2�J��R,#D��j���Č A��ĈS� 	�D�EP�<��y��}���nI�л����
9e��]ۀ|��l6�X}�|�l��N%
f&b����?C�x���s����]��`�[� �� r�-@�Ur��l���:@کzy�@�(9�rO���v����A[��7,�;��X_���Zn�.%�K���nl�{�2�!�����r��\ �� �^� �{���\�g���)a����� {�?���\���/up�ˉ�1Mr`��SUa���s�*w��6��j��w�l'��Ą�\^\�ٙ�33$�M�xGeMcz��<�T�������\\O/6:�[�`|��0�v���:ݱ�k-Qգ��f�\a.�✴M�ҥ����Ee�e㣤�`�;� >�ݸ϶���d��_�in������ĒQa�M��<�`w���g;�i������>]k�{�b�>B���͋ �[�`z�*�U ��@�`���?��|���< ��ά5|��q)�f��{�2�A*�ѲZ�ݝ׀���O�V����ܓ�{��� ����e$V I%Hąd�aP���W4&�#17�>�8�a�A�0��1bs��Ѹ�v0����JT1*��0�Fl�aVX�!1`E�����ӧ!eH��
T(���bh c0c 4���"���z�0`F ���H2��$�,���s|6|�B:BR�CA�����y�qt(Ba�W����y�M��K�`+#��7�6pͫ���Bx�	䌁�1$\T d �H$��!=C����J���	T��?X;�66��=&-�հ         �$ְ  M�f��Y�vZyᨮܶ'��z���Y��X%ʼ�D���٫mRy�nր�  ��     �      5���Ye��u퀵�t�;:Q�/�^k�g-ح�Z��[�1����D�oJYn�\\s����K�cr����]<O�[ˊ�c ����;Z�62��n�!VvOFĠ�����o[9��ۑ�h�Tnp�Vn�N�D�ƹ��qz�lvĖM6�I� 6�����q�]�;�wWlT�4@E�۹6�8��YrlYN�wbcm]i���;���nt�r��t���Z(n{6�4���n�����L�5hKF�-�|��W��V��]�uӂ��pvj���u�;��ݣ=�;�\'Y�"@)��@�UK� l��lN���{\�.���c
�� ڠ����s=bݱ��蹪�ʛ5@c�G@2�`��7(Y �7J�����gf�D�fJ�9�ܙ�B��q/�%�ٱ%E���ջ-�U��B��v�5�کʷ<�K/;l�u��b���lv0�Y��V��t �c�����tZw�G@br���n���.jZ�gZ��l�+UJ�յY���2�뛫$u�oN�{86Ͱ   I�K6���n��-�&�T�̓Į0���Q�t��-��&m�.""R�����D��u5���W�=�9�!&cL��AΎ.��ĞXݳІ�u��жk�6�l�uՊ^Nk��;FV�k��\ݎ���S�Sq��䝫4n���T�)y4"p�2 :�팮
(u�����y�:�lo�A<��UJ
7^�q����9���:��v�)�Ѱ�`;v�t�j6���]���.7.CX�vѩ��qv�g�1����;qvBdG9/i$�s���Xl/5�������� 8  
]��&��D֦���Љ����J)�&  � �"���8�О
x���U���)��w��w��ߩ���t˛ A�̖��Tδ�1 UX˭0�Z;�ˍ�e���[��I�z�62�b.�H���b�q�笳����:���g7aM���gB�n6A+2�j�@]	o�t�c<����]�Ҝb����%>�t��,3�����<Z0w*����j�ڨ�sf����gvĂu�L�Ύ��wF�Fـ+�2&3V<��L�R�[7{���w��]O%lk��d�G<l��e�Y���H^W7J'(pؠ��$OfF��V�嚇�%��� ^�v��\�u��?/�B\]�y9�`��6E1R�����݀|�� ��f@=Ϫ�{:��)q.o>G9�T~��S5%T�������j���,��:��n��É�E�REr(�*iX|�7���IVo��,�U�~�u`~ͅ9#�L@��i���qv }���[2����&q3��^���ܵ��R����\���Z��ۻ7g��u��B�g�]���{�pIg����H�u2�)nq~8��bX��_�]�"X�%����"X�%�����iȖ%�b_}��b���-����"�+rT �y���ı,O=�xm9
�ѵHZ��ӌq�1HB$a�j�K��3�ꉡD@��X�br%���s��9ı,K��O�m9ı,O>�z�㉜L�g���IL���F��r%�bX����v��bX�%�ߎ�iȖ ?� dL��u���r%�bX�����"X�%��{:sSY2SVf�n�sWiȖ%�b_}��bX�'�k��ND�,K�{�ND�,Kߵ�nӑ,KĿ|I�N�2�ђ�upֶ��bX�'��{�ND�,K $��=�����,K������Kı/��w[ND�,Fqj�y�#���)b��2�ԕK�;��mn.�2�L���ӷa�mm�;Z3sZ�m9ı,O=�xm9ı,O~�}�ND�,K���u�_�AB(�&D�,O{�߮ӑ,K�����2���K��[.�m9ı,O~�}�ND�,K���u��Kı<�]��r%�bX�{���r%�bS�}��A�X������&q8��~;��"X�%����nӑ,v(l<Q"рUD�@$;���\4�AJ)UhA�_?A`�A 蚉��~��Kı;����r%�bX��:w:�3.e�f��ѭm9ĳ�U�����Kı=���ND�,K߾�fӑ,K�H�B$>���m9ı,N����Y.$չ�$��ӑ,K�����ӑ,K���ٴ�Kı/��w[ND�,Kϵ�ݧ"X�%�����uL֤�a�����Ý��j�E&We;]tJ[���k���27 ���z�����~oq�ı=���m9ı,K��ӑ,K���w�i� �
�a�L�bX�����"X�%������k%�!�d�q|q3��L�}�\��Kı<�]��r%�bX�{���r%�bX����6���*D_��`!���b_߉?d��e��,�WkiȖ%�b}�_��iȖ%�by�{�iȖ%�b{����r%�bX��~^�����&q3����x�Iaj�7n�v��bX+�"ĊdO~���iȖ%�b}����r%�bX��~;��"X��
x�f�k�w�iȖ%�bw��\�冤˧5-�Z6��bX�'�}�ͧ"X�%�}���r%�bX�}���9ı,O=�xm9ĳ��_�������A���[��v�i�;6�ؤ:�x�5�%�Z�K��T�˲������������>6K �v�8�q3��L�~���[ND�,Kϵ�ݧ"X�%����"X�%���o�iȖ%�b_C���a#��������g8����w�i�������'�����Kı;����ӑ,Kľ���m9�&q3�b���"�+rT �y��%�by�{�iȖ%�b{����r%�bX��~;��"X�%����nӑ,K�����3,�D�Z���ND�,�ȟ~�?M�"X�%�}����r%�bX�{���9ı,O���6��bX�'��t浐��jk	n�����Kı/����r%�bX�{���9ı,O���6��bX�'��}�ND�,K�ثF%���E D"%
�ޗ��~M��n�0 :t����v�m�6��m� ќ��;f�xӊu�v9�ӷN�/]����qY�5J:tct�/b0qm�^t�&�;���X�ݹ�=l�B"L͞u݁z�϶�%��^y\�����<����Lm�{x��OgB�E�@p��d���]���Bq��+jI�:Q.�EM���fݎ�rjwb݋F���,���
M���w���i ت�~X��) �%�$����䃑ϐ۬�G
� ����l;j�h��c��\��+��#۵�2�v�3u�k!m���q>�bX�'~���ND�,K�~��"X�%��~�f��@�DȖ%�}����r%�bX����?�j;T��%�/�&q3��[� ��r&D�>����ND�,K����m9ı,O��y��Kı=��#�T��::IVq|q3��L��~�fӑ,Kľw��ӑ,h�lS�eqX���6���q6���"&Y&B�i7�_�a�L�����r%�bX����m9ı,O���6��bX�L������r%�bX��>;��&e̺�ԓZֶ��bX�'����r%�bX��G�����,K���w�m9ı,K�{�m9ı,K�����V�ٙ��k�l��r��3��ҥ�&n'W��C�*��q�j�]�vݚ�r%�bX�}�xm9ı,O{��6��bX�%��bX�'�����8���/�瞒(�Cv�Ij��Kı=����r����T:�#�_��O"X�������bX�'����iȖ%�b}�{�iȖ%�g�Ǘ��6���n�)�_L�g���[ND�,K�u�ݧ"X~a�2'{���"X�%������r%�bX��:gr��m�Y��ӑ,K���w�iȖ%�b{�{�iȖ%�b{߷ٴ�Kı/�w��r#8���&�ǃ�5��D춼���,K߾��"X�%���#�����yı,K�~�ӑ,K���w�iȖ%�b����-�Y�f��]MZ
0��z��٬m���'�����~�zቺ�q��XZH�X��ttr��]8���&p����M�"X�%�}���ӑ,K���w�a��<��,K����iȖ%�b~��M��Y��f�&�u�M�"X�%�~���Ӑ� @ ș������9ı,O����ӑ,K���o�8�8���&qv#V�q���`�۴�Kı>�]��r%�bX�����r%����Kl2�~"N��?�CȞ�߼���r%�bX�����8�8���&ql^��UnJ�<ֳiȖ%�£"}���ND�,K��o��r%�bX��{�m9İ? 2'u����r%�bX�����\�Y��n�)u�ND�,K��}�ND�,K�.}����yı,N��߳iȖ%�b{�{�iȖ%�g�}�q��U��Y%��T�9l��=�u'd�vl�qZ�%�yc���B�;TTa-ֳ56��bX�%���[ND�,K��{�ND�,K�~��"X�%��{�ͧ"X�%�}���w!m�˦۬��m9ı,O���m9���� 5Q,N����ӑ,K�������Kı=�{��r%�bX�o��j;T��%�����&q3����ND�,K��}�ND�O��DQr&D�>��6��bX�'s��ٜ_L�g8�wČ_1J��vIM�"X�%��{�ͧ"X�%��{��ӑ,K��;��ӑ,K��	�@I:�U� �"k��Ŝ_L�g8�����0VFJ�(���ND�,K���ͧ"X�%�$����m<�bX�'�~��iȖ%�b}��iȖ%�b_~���Z+aq/,��0��a�}��{v�\�\��Ӻ�v#����c���٧iȖ%�b}��siȖ%�b{�{�iȖ%�b}��a���&D�,O��߳iȖ%�bw�Oں.$շBf��ND�,K�{�NC�@?�*$��j%�����iȖ%�bw;���ND�,K��{�ND���&qw�G�Z4�8�8��%��߷�m9ı,Os��6��bX�'���6��bX�'���6��g8�����>�QҺX�풙���İ_� ���}��m9ı,N��߳iȖ%�b{�{�iȖ%�b}��iȖ%�b_=$��[u2��35�ND�,K��{�ND�,K�  ���@�{���M��,K�������Kı=�{��r%�bY��{������������0l�E1�c���v�V��b���Sg�bg�pj�[��!��������N�75,��-�n����Ʊ�,<]����r�X��;2��l֮�����#Ӣ|�.;���nz����:�!Z���J�&�������g���G ����_=���Cqz7An�q�.=�l�n��&���wognz�-��UV��ow~�����[����lt0Z�+�a�yŻyW;V���Ӂѓ<�v{uW�]�9'W)u���,K���~��Kı>�۴�Kı=�{��r%�bX�g{�_L�g8�wČ_1J��vLѴ�Kı>�۴�?	���H�&�X���fӑ,K�����ٴ�Kı=����r%�bX���zG;UD�8�8���&q~�{��r%�bX�g{��r%����>���m9ı,N����iȖ%�by���:�3-�t�5��r%�`��02'u����r%�bX�}��6��bX�'��{v��bX�'��}3�㉜L�g����A[qQZͧ"X�%��w�ӑ,K���o���%�bX��]�v��bX����zg�8���.���Y,���ѓ��nx��05�0�q��c9�u����q�Y35�����5w̹0��jR�q<�bX�'k���Kı<�]��r%�bX�g{��"șı>�p�r%�bX�����B]]]Ma-֮j�9ı,O>�{v��A�(�c�5��;��ӑ,K����iȖ%�b}�w�iȇ�L��,K�ğ�����e�mֵ��ND�,K�����r%�bX���xm9ı,O����9ı,O>�{v��bX�%>����Gajpv�fq|q3���.pI1@u��zm9ı,O�����ND�,Kϵ�ݧ"X�%��w�ͧ"���&q~�����)Y\R��*�/��,K�뽻ND�,Kϵ�ݧ"X�%��w�ͧ"X�%�����'8���/�}�zҹ+r�;$�;�y���n"7V�7aHyAT%P�X��K8�rB\I$����	L��8�+c%�Q;*�����X�'{�߮ӑ,K��;��ӑ,K�����"X�%��{�ND�,K�'���ən[�R˭]�"X�%��w�ͧ"X�%��~��"X�%��{�ND�,K�u�ݧ"� �*dK�}�~ֲ\4I�n��k6��bX�'߻��ӑ,K�����"X�p Ba��+�,*B��
�1�jJD�)f
E�!�ޚ�C�D��7�CC7v��� �!!BB�#�2`V ����0�<�����qvh5˽�8��	%�H$�4q�����6��AH�9�	P��w��60I$C����a8+�<6����801c�!P�%XVT%#P�aA��H����ʞ:!g-���EL!�����A��J���ʑ��=O!���3U�HHiN.�ie�2�:0�iB��z�Α�U�*�P1႔@����=�SJ	Tة�� E��A�b��@
��|<�y��>����Kı<Ͼ�m9ı,N�۾�3	0�-֥.kFӑ,K�����"X�%����nӑ,K��;��ӑ,K���I�?}���ӑ,Jq3����_[�+��n�j�/�&q8�'sﻛND�,K�c�~��6�D�,K�߷�m9ı,O����r#8���/����F���n�Pm�Ez[���qX3�ێ�ܻV����k [27�3Y$��e�m��k8�D�,K�����r%�bX�����r%�bX�w��?��DȖ%��;�ٴ�K�L�k���O�!%R� �����g���fӐ�9"X�����"X�%��;�ٴ�Kı>�����Kı<�������3R�sSiȖ%�b}���ӑ,K��}�siȖ��2&D�~��6��bX��׷��~8�⃊,��1 ��	�$�.�Fӑ,K��}�siȖ%�b}��siȖ%�bw��iȖ%����Z/��D��߆ӑ,K��	ӹ�ən[�Rۭfӑ,K��;��ӑ,K��� G�߹�m<�bX�'~��iȖ%�bw>���_L�g8���@��P8U\U�S��a䳃��t�y�3�G:�2��W��n�ak��PV�TD�g�8���/{��m9ı,O����r%�bX��_v�9ı,O���m9ı,N�w�j��F��/�&q3��[���ӑC�G"dK�u��iȖ%�bw?~��ND�,K��}�ND�,�g�o�������7l�g�8��'~�ݻND�,K��{�ND��DHdL��o��r%�bX�����'8���'���n��6岼��K��,S� j'��fӑ,K������ӑ,K�����"X�%��}�siȖ%�bS�����s4f�fK�fk6��bX�'�w}�ND�,K�c�߿xm<�bX�'���ͧ"X�%��w�ͧ"X�%��ٲ4H����=���ӽ��?�ۗf��Yq�.Qև� t�vͪɍ��j��'lg�L�g�9�ݼT�v2�vV1��>�-��;ԛqۢ�v��>u���J`�����Lj���|����I��+m�^������ƨrsٹ\�sՈ�8�r�H�\:����۝��Y��1�:�$A�nÀM�8�8y�����X
��c��/�q��u*��^��{���w��������F�M+�ۣۗs�eѬ�M�%��F�-s��{8s��������7�M߄3Z��Ԥ����%�bX�~���"X�%�����iȖ%�b}��siȖ%�by�wٴ�Kı;�f�r�����Vq|q3��L�����/��)��,N��߳iȖ%�b{���6��bX�'��xm9�`@ʙ������.Y��Զ�Y��Kı;��~ͧ"X�%����fӑ,K�����"X�%��}�siȖ%�g�����L����l�/�&q3����fӑ,K�����"X�%��}��ӑ,K��L��~��6��L�g8����t��j��H�q|%�bX�w]��r%�bX�g��m9ı,O���m9ı,O{��m98���&qvn��(�Q��J5r��U��lt����U��H卮)"{27b��!b���㉜L�g���p�Kı>�����Kı=�wٰ��H�ؚ�bX�����v��bX�%��'�?�Im�˦ۙ�k6��bX�'���6��T�$F,R!� �&D�>��|�ND�,K��~��Kı>ϻ��r%�bX�����##�Z��Y�_L�g8���iȖ%�b}���ӑ,�"�!����?fӑ,K�����ٴ��g8����Č_1KI�c��.D�,K���6��bX�'s��6��bX�'���6��bX�'~��6�L�g8����v�����Kı;�w���Kİ� �������{ı,O�����ND�,K���6��bX�'~�s%;.i�]+�9��M�N���^�۵ۻgz5�IuKrKh9v[����L�� �����"X�'���6��bX�'~��6��bX�'{���O"dK���~�v��&q3��_�o��]QJ�[qQىȖ%�bw��iȂ��@2&D�;���ND�,K�u���r%�b�ų���/�&q3��^�wΖэT[�I��M�"X�%����6��bX�'~�{v��c�Y�F[Fؤ �ls�<������6��bX�'������&q3����}d-!b��h�r%�b"�2'�w���r%�bX��߿fӑ,K����fӑ,K�����"X�%�~�O��Kl��t�s5�fӑ,K��;��ӑ,K����fӑ,K�����"X�%�ߵ�ݧ"X�%����N��*��hM������wȥ�Vm� �:�u�6v�*�&�&��	&L�\׈��|��˙U,R�,�-8���&q�����g�X�%����6��bX�'~�{v��bX�'s��m9ı,O}�fe�,3Z��Զ\��r%�bX�w���Kı;��۴�Kı>�����Kı;�wٴ�_�ș����ٔ��&]d�P��6��bX�'�����Kı>�����Kı;�wٴ�Kı>�{�iȖ%�b{���팹f[�R˚�ND�,�02'u����r%�bX����ӑ,K��{�ND�,.�O��S�8���3T�R�E�BP҂H|1���4��������O߿w۴�Kı?a�guta��շBf��ND�,K�w��r%�bX
?�������,K���~�v��bX�'s��m9ı,O;�?�5��k'��Q�v�+���X�i�s�r1n�ns�L�:�P�^�-$��w�%�bX�w���Kı;��۴�Kı>�����I�L�bX����6��bX�'����k	��S&���Z6��bX�'~�{v����G"dK�~��6��bX�'���ͧ"X�%��{�ND��$���|v�$�1��f�pI���͉ �'����p�X��w���6��bX�'����|q3��L�k|?z7#%R� ��ND�,_��O���ͧ"X�%��߿p�r%�bX��]��r%�bX�g{��r%�bX�����Xf�3�m��ӑ,K�����"X�%��뽻ND�,K��{�ND�,K��y��Kı.���
�Ͻ�߉�\� ��]5�i.V�"���	  K)�.�N�SZyƝ�V^Ѡ3�����K�-��]	j��rv8��zSt`m��^Gcu�umݷl���S/Es[�XwcV����<\l\v"]e��u�C�U�D�7Z�b�*6���>��#�EmlM;=9�0ggb��v�Z酮gk��=��Kv+c��휝�׆ۍ�m.\$�T)������;"���*vuƶ�U��GJ���sZ����$Sz��2d��̚�&�s4m=�bX�'���]�"X�%��w�ͧ"X�%���}�ND�,K���6��bX�'�N���˖e�u,����Kı>�����Kı;��iȖ%�b}���ӑ,K��u�ݧ"X�%���wWF4�ۆ�3Zͧ"X�%���}�ND�,K���6��c� �.�j'�����ӑ,K�����ٴ�Kı;��H���A[)�_L�g�%�q@ȝ����ӑ,K���_�]�"X�%��w�ͧ"X�%���}�ND�)��/��)��Q�R�7l�g�8�K��{v��bX�(� D;�߿f�Ȗ%�b~���ӑ,K�����"X�%���v��r�	nI�es3���\��n�`�����Mj�7 �	�� �[N���K�,�����7�����{�ND�,K��}�ND�,K���6�<��,K�~���r%��&q5����J��A�%�����%����ͧ!�Z�U��@� �lO"X����ND�,K��fӑ,K��;��ӑ,K����fXr�4k0�Ke�M�"X�%��{�ND�,K���ͧ"X�,2&D�~��6��bX�'�o��r)�L�g��=#�ND�8�8X�~R*���O�����ND�,K�fӑ,K���fӑ,K�����"X�%���s�2�n�In���"X�%��w�ͧ"X�%��{�ͧ"X�%��{�ND�,K�ﻭ�"X�%�|��;�kSF�fr�f��0{e����6���x�����qn�P�Xce�\�@=n�?{�7��bX�����r%�bX�w���Kı/~���(����Q,K�fӑ,K������&��eԒ�jCZ�M�"X�%��{�ND�,K��w[ND�,K��{�ND�,K��}�ND�,K���9�2�Z˩��Z�h�r%�bX�����r%�bX�g{��r%������2��~"��j&D� *f��4+�0��X�����7�=���r%�bX��w��ӑ,KĿ}'�;�-�S.�m�f���Kı>�����Kı;�wٴ�Kı>�{�iȖ%�b_n���8���&���A�)T�H=k3Y��Kı;�wٴ�Kİ������O"X�%�w����Kı>�����Kı? 	߿~���i�:-���\�mu�����Rv��7K��f-��ziue5��������yı,N����ӑ,KĽ���ӑ,K��;��ӑ,K���g����g8���j�H�S��Q9�6��bX�%���9"X��߿fӑ,K������r%�bX�w���O��ș������2�n�Iu�kiȖ%�bw?~��ND�,K�}�ͧ"X�%��{�ND�,K�ﻭ�"X�%���wWF4�ۆ�3Zͧ"X�%��{�ͧ"X�%��{�ND�,K�ﻭ�"X�����Q�b���}���&q3�ݻ��c�7h)e3��%�b}���ӑ,KĽ���iȖ%�b}��siȖ%�by��iÉ�L�g�}�q�Z�#*�K%h-��&��b4RvI�Wm	��:gˤ���e���(�6햬���g8���w�iȖ%�b}��siȖ%�by��iȖ%�b}���ӑ,KĽ�O��aH�nYnq|q3��L���zm9lK���fӑ,K�����"X�%�~���iȖ%�bS�}�R� �����g8�����fӑ,K�����"X�B"_�w����bX�'s��ٴ�Kĳ�w|HφԪȥnS8�8���s�D��߼6��bX�%��kiȖ%�b}��siȖ%�b}�wٴ�K�&q{ڳ�9���`NJ��㉜LK�߻��"X�%��w�ͧ"X�%����fӑ,K�����"X�%���xw�\XhIg�!1 Fzލ�A �&��,�bk���b�9��bF$�~�d���#�6���l�� 70$H�!2��1*h��<:��U���i�!����\�"����1&M���%,J�	����c���`۷�hV�@         m%�  n�֑b��:��1s��ݦ�[H\��� ��!�qvDr2�����۳ �  ݶְ  �  �     �`�t������H�lU���5����s�q`�V�h�۱�6�v�ٝ��Dvx�V톥t�ݬ=a�+vH^�{�ҁ��4�5AS�`��&�l�l؝\����W]Q5��<i���`���\�v�v�{<a�չɜi�&��N�.��R��"�jMt�<��z��T��`h�m-����N���I�IŚ�X��4�Rr���q�=�ۣǷoi�(�f%�#\]d��cu�'��C�&�[4���V�wAv�Ӥ�|�s���3ͳ.L�b�vCѧŝu�.�}�Z�:n�4��oM���ا����뜥�som����"f@7'%���jW�^k�����+���n�,s5e@v�V��vP�۰9�B�{6�F6���jg1����ų�]@r���7mv(���$ʖ+��נJ���'diGc�P�{"��0�ֳ嘤.j�����"�\����e�!wn�t�zӅ�ɥ���n�]n��ez�v㎀��[l츶�V��v(���̜Ma��;�qQ-P
j��.��UT�R��U�E������p���T�l   m���m�۶d˓�@�U����<C��m��m�PvN42�X�nͻg�X�6[j��ӽѮEM&n-��,d��S��]±c��u�I@���1ۧ\�ε֋�k�Vݲ�#�\n�5�+�rq���*�pI��pRY�qV;j�9l��iЎ@�۝���lv�R˃��Y�0��ym��)K$�n�q,��ҕ��IeY�*]��4���ؽb�uZ�+�q����jj
� R�v]��6�Σ	�.��v�杖IZ3GSZӴ�I�m��-��   ��dut #>�w��U�D"��` ��
�M�
(��'�m @<�{���P :j�6����YU+m�H6����Z[���V���g��V��UЃ+h0����T6A��]@.�խ�ǳ���n����b�c�`���li�͒�My'�v���)���Q��[�8u��x�瘧`]pV���8Z�X|;s�n�A��q�fu���;���L�О�kv��K�s��礉oS���k3333T�ԙ�ED�'5����8��^��y�gAv�A϶u \�q.��VH��(@$m����!z�5~ND�,K����ӑ,K����iȖ%�b}����?��L�bX������"X�%��>�?j��&�[p�&kY��Kı>����r%�bX�w���Kı/����r%�bX�g{��r'� eL�b{����ֵ$��2打Y���Kı;���ND�,K�߻��"X-�b}��siȖ%�b}�wٴ�Kı<��3��u�]L-��kFӑ,Kľ���iȖ%�b}��siȖ%�b}�wٴ�Kı>�{�iȖ%�b^�܅�ԙ�[u��m9ı,O���m9ı,O���6��bX�'��xm9ı,K�~�bX�'~��e3;��^��sj$8z�\63����ռ$݁�>���#p���U�w}���~8����1��"X�%�߿o��r%�bX�w���Kı/���� 
O"dK���~�v��bX�'{��弖��e�]J[��ND�,K���6����!!�-��BZ�(�"����Z2F,����T�?
x�'�,K��9��"X�%�����iȖ%�b}�wٴ��ʙ�����f\e�rk$���Ѵ�Kı/߻�[ND�,K�뽻ND�,K�{�ͧ"X�%��{�ND�,K�P�<�0��m�����&q3��뽻ND�,K�{�ͧ"X�%��{�ND�,K�߻��"X�%��wǫ�(^V�TQ��{�� ��K7w��sj��6���|�*&��j���h�m����rf�;�*�!�V�8n�7v�79J���[@vr�S ����v���봀}z��ǯjh�ST��ίW��2dn�����<۵s�D&��$��	�R[�k��0�ۦ��BG<3���@�Z-
�}��f����nI=�_vH�V���Y���o�����X}�VĹ���ˊ����7w�&!\�Z-��ِ��`�� ��t�?����=i\��b�Q����P<��Cl�p�,���nr����<�W6�S�`�`NJ� ��׻� ����8��]��ݵ`nJ#g`�1\��*���6���A����y�j��{�0��M���ycqQـ}�t�<۵fqqD8o&�q��`~��ĕ4T�����a�9ľINn�U����`{~��ܛSB�'�}���~�uL�
;k�Lv�V����:�� �ݤ�� ��5��@�ݐs]a��܏7%���ۄ��3l��Bjf�W [K���,7B^��0�ݘ�:e��ݭ�Z�� �3f�3L��)����K0��L��� ����9[\�Q4��=�x��OH�v�Ǽ��K�j��F�́������#�,*��rU�~}���[���2���%�3?+2Q9�o�5-� �mp�� m� ��߳rM�jT��K@�
���b6VRA���$$��"I2BJ *�F7�� X�L�@�,��DY$�R,�a!�0$%5�(s���� �@cs6�r�W�H ����EZ(yP��AX�m,q�z���(P�<�am��F�u��csn%�ΏQ-�
�m܍��X���f�
3�b��*�*.��3���[c��	�Q���:�Z ��🏪�&�[@k��u��^�z�8�������<��)\��e�w+^^K��6%��q���`���݀l�w��������{�~;s]���u�����^�:k�ω���=\逹'�j�p��������~}�"�պBU����_�v�Ǽ���6���T�z�1=�� m� �{�lCnl�t����A�x��P��JD�k�`{��^��?ˉ��ٵ����j�:��#�E"k��4����]��� ]���z\��f�R�2ET�M��Ι`j�՛���7'v,Cnl���TT��������n����$n(�s�ݗ��4U�`���ݜ��r�7[jU"�Q��0��,�@9[\��@-����bf�I�\��}�}��E�	�����)kH��uj �� (I	�0��F�tK�PQɨ�ĸ��2;����e2��n����&�6v0�"�j,�ݛ��0�&���,�=�u��muNK��0{�z� m� ��PV� �Ӻ�e�Aʄ���ŀ�?ۗ�#wf�~t���H�T�PA@�9�a4��35O4t�mgj�ғ������"X�Qʭ�
;T�k�`ٺ���z� m� =��������{�������ِ�n/W6d1i��eLR�T�b
���{�_�����7)'�T�Ġ88.u!@�����.�^��l��ojXH��)��%Ǿ��V9̋�ۛ��,�����AR
&iX��Xq}����76��;���������r���J�N�:�]�9D�0����ݐɮlZ�4���r��e� GyGd��5�ޘ��0��/qs����=�k]��ꜗ�9
"j��m�/�������T��Ł�������\,�;9P���?w�ذ�j�uv��i �^���kX��UER�����6��m�,>�Ĺ)T(�T�;��7$�:|g섶�'���{����ݤ�� f��?�8�o�����b��*�����}
]uf1Y�7֬�Yj�vn���L)ۜ�=e�2�*IT�b
���������ݫ�j�r��z�&��=c`�HOKͻW���7gv,�ݛ�L�7z���G �rU�n�׀u��[v��̀^xV�0`���*f���6��m�,6�Xo8�2�# 4��T墱�Q7+�7v�~~v�帰=�n,�'-�$�����Q��vmt��8$ ���6�ؽ.i$6���Z��>ﯝ�t݁����I.�˓�L�H� ݲm��gTLIZE��֐��d΄�m���`�s'Xnz�<����l�&m3ϳʑ�S՝᳎�T�'XF���;�ۧ�ז���Mk��t�GF��]�kkD�X��Ѱ]��خ8��qR�{��^�Z�_�{�������s[Y���j�;ԧp��j��9��J���L�sT��uڸY@vr�Y)�o���`�u��j�[v��z��0�i������ܷ�9���Ł������j���Z����9xG����<m�@=z̀Z�P��to�oBf ����t���Հܷ$�ӎ�b�Ǧ�LX)���"��&���d�j�w��m�@/Z؜Okaũѫ�˪K�dzK����j��wE#7A���a��Y���:絸[��~��@;�� �� �f@/<+u���������	!"q$���*��9���\��}��ٹ'�g�]�*������X�(��������s �T��P��3^����L�`u�ڰ����e���|�wi�y�{�[b�X�*c�ڰٺ����fG�32��:��X�s*&��YFgu��r�]�h�ISn���P����2I������wd#7�#G�o��U@-�H�Y�]� vS���UIBF�-� �ۦ��;��,ޞ��;�n���8ٽ����RK+�h���=�-X�qe��$q� �
�HV��!$aRVW|=��=>�!�hK=瞍�
f�jK�m ��" �l�J�dM�>��L���/��S4!))(�9�(8�5����� ���d1\����
��+(���
� �+
��0 D�͛.�~���0�#1�B"��� H����C��ѧJE����X�� ���oa�	|��!q��S�f��&��m��A�$$�a2I	$@C�_� �T�W�h�*�����PڻUM"�
�Q�)�����
���S�T0M*�����n�I�~�� ��#�,*��rU�n�׀w��X�e��/����7%3� �������@;�� �� �f@7f��?ˋ�'��=Z�����H�.���e���K�]0�qu����39�Ŗ6�V�tW��
&��z��?ow�7^��u��w\�P��h'e_���s�rwb��;�`?:e�����lY�L�Bz�ryڠ�j�^�H�Y���̬bC��M=� �;T��@=ź�s~���9���>��}��~��S5$�D�5U�X%�.{~_��9�`{��X��c���һG,C�����"��WQAEi�QU�s�Ȳ!3U��=4��%�+1a�=>�����j�w��z� �Wds���P+NJ���y�����)��Ł������j�nP�a�!<��-oT��P�i ��2yڠ�Y�����6i�=P�i`u�ڰ���ĸ��w��ͩ��=m�n�-z@=z̀^v�{>��I��k�& �o��+m_~�����. Ӡ�V�]�p�,m�	� �\�pՃ��n��%V��̽W�eӃjn�
��a:�`k�@gj1�]�/J�/�,G%s���%�W $���{y���h;GAg!�a^�n2��/���g�~���v��9��@-�)�G�`��2Y��j���kE����S��n�!�ô�T;cu��ꕥY�u=���{w{���E�ѓ]+4q��8�A���T-q0�h�LA���p�UuO'Yrջ���@;�� �v�^� ���l/u�^��u��L�:��X��_��_L��ژ�341MUE�������j�~����;T�J�P1��V�a�= �f@/;T��P�i �ski�5�%)
�4��n,�s�_s���s��G��~����Ձ�9	��*�����%��m��I�ɮ-W:����b]r��P� ��"$�$����_�og���X~v�s�~��9�`=���S��MB��ܓ�~��z��:PQ.�."�ee�2}�`{��_�.}�ɓ\���4S3U��,����m��\\M�g��o���{�� ��Lr�V�I�o������ۦ��d �v.���O&�=� �:���.%�8�7���m��[��ӓ��&����Zw2p�N����ⷆR�:붮n\���%n.٤yI���MUE���_���[�����̌{��ǀ��UX�[��?ow{��"s���E�ۦ^s�_s���G����`�T
Ӓ�������;�n���"�A��(]���3ڭ��� ��s���EL�X|��?VdX�XX~v�1$�ğ�}���M֯#rM��n�`?yڰ���}�����.$���6�Y��k��:٫p�6���75C�1P���l�r�N@���I/���>�ډd���U5K�}����n,�n>Iq%�{�ŀk��[b�R8T�k�`]�|�Pm� ��d ��]������:� ��u�����s���73mX���Φ%L�MSU�m� �̀Z�Pa��������&�cM�@/u� �ڠ�� �ِ�뻦�oRg�+��]V\�� ��"�񵳛��6:ۊ7��!/�������8Z8U�IW�7gv,�n,۵`?yڰ�f`�C[�E��_;T�f@/u� �ڠZ����$��Ğ��̀^�2k�@*��^:���&�f�ST�7�Z�ww��ݝذ5����.?{��`���� ��M�^�@-v�V� �ِm� y������~N\ h��l���^D`��T�UQ�@�+C"�K���v��N;N��;��ݺv���`���[S�'<]��,#�q���%lL��M�U+Z�.�:���`W��C�ۍ��;&���{[�WlPa�Q}�^�MzDR�%���i)��pX�ngllY����g�ϫ�?n{=&Km���՟bp�vhg�"�6�,�ݲny��k��UcV������h䭍a�A�]XHy����Qu��	�\��4�͵]l��u�ӹe�LTMTt�y6mڰn���d7gv,5mLJ���&"�f��m�Pm� �ڠ[\�J�Y?4��lXh�rm� �T�k�]�ŀn�]��Z�$� ݛ��pۛ��Xj\[;��V�fcs���-oT�k�[l����7f��>��j�KP8Ud+��^
���n�鮧�g�uJ�s��9�q�;��nm�7���$�����̀[l��u��v`��m��H�h+-XI��}�؄Q�S��qrx��.-�?l�Ł���`6ݫ�z��,�&n$�^�@-v�V� �ِm� ;;b�F�{�5�UE��6mڰnՆ��xX�������%���,vِn�U��.[��n�Ԛ7Z�H��������s��sR[s�%��u�`�r����rJ��:;V��� �� []ϐ[w4{6���X����܀w>4]�8�ِ�ڿ�ų'�&7�30LW(������?f���ng�"��O�D9ϼ�1`ݺ`��u��j���`�v���X����Ĕd�6�M����1�
Հowq`ۻ�>��=0�w�Ӯmj;A�q5�vK�$�X�2�6B��]�un�#ج��3ıʣ���Tn�Հw��`ZW ��� �l������f�TX��q�e���t���)���B���j�~n՘�����yZX�́��kq��rZEr�V��ŀw�n��}~>�7$�"�@� �o��^��{گ��E��V�	*�;ݴ�Ur� ��� �ِ/s~K���]��қ"�sDkA���9����/N�.��c�[A��n��ݔ2^���Ḿ��ڰn��/��Ȱ2�y��j��[0�w������W-p
�[����ؐ�C�rm� Ϫ�Ur� ��2���E�Q�T�V���<#ɰ?6�Xj�f<���jr���P��Mn��Us��}m� ����=�=��I�)�X@!���5IE�"A� ��i I@���d0`� �� [��#	�<ԃ��Č �1�v�0b��"@�Pڒ��K.!�&�PڢRA\d�\�BAH#���Be%G
�hI�H���'D*R�dp �FR��o��|�I0��kV���U�.+          m���  �I��5h����U��^���,y��H:v��vLeU5�4��m  ��  ��  ��     D�`���j�׬�֑�\����u��L����sCX�Ep&���|�7��ӹ��M�멇!s\q5����QQ0Q�zq�J鹭��ntxm�`V��`�v��%;�i��w����ܪ�cO7�W��T!�9v����1
ɚc���X����/6Yx ���"6��p�ِ�*8*퐠R�q�c�ï��:��;K}-��1yIo]$�@�lh�c��&ye|J�Y�"Rth:������^^�w[���A�*={!��V��$ �kuG�H��e�f�s/޻]HV�mp��H������n�n�??}+-�L��6 �>qo>�5
�^s�r\����%i	�QҲ]�n{a̸�F����lCKE5�a�S'f�-��� �O��E�R��l
��VzR��D�-痛;��nQ�tc�ptgu7.؎�͇��I�u-ڲq��7J�O^8^���l����p�9�,^CgS;\8�G������հݳP�g�� ��ɺ˹٭�p�N�ٰk�q$�C��V���Q��3��kf�]�}��o�  KW�CAڗd�{j�U�{��KW^M��nܥè �c�A-��4�%��&;lr�b]�[�'h���m�E�q���8�t��$Z�S��X,�h؏P����c��7n��4����l`�.���OU��/��O\�quV
�؁���5�Q�5�rN�<x�@h�m%��wl��Uq�T�{3�-��+���y3�q�:�=<۰El��v��rm��Z��4�ʇg��7 �[�����������Y=]��)1�j�]�H-���   �8�I+k�9�8
����E1T��� z��xuJ�'p@��PR�� ��D0>С����2� �a�ՔQaK� �u�m\t�=�anN.�k�*8��u�h�H�9�p�n�x��Q��O�-����\&"']��� [�9��s�<]���Vk��L��a�9˵�^'�{b��5���q G��Z�U���{(Uۮ͊1� �sˍݜ�vɌ��{/nl񸓎ћ�v��|p�X�ݐ��Y�kY��Z35�蠜3��^��v�7O'=�|}��]lVY�s����f�r���ɰ�v�c���Sm׏_�������f@;�U ��W ��Mn5��KH�NY*�7{���ē��yF'�`~mڰ�3¤�7�{���@*���>�̀[�d��ͫ�1����u@*����v���Xb���Xy�J*5xۊV���ۻ� �.s����|�vo��Wv`?��KB��id7U��dw�^��F�].S�8�$N",��L�e��%�ڭ�lv���`��X{:��pל�\_�;����9�UL��I����� �}Tx�Uή�l��wy% wǔ�VF�d��;m� �՛6��j�o�Ձ�ϜX�tX�-z��x��>�f@-�2�Ӻ�z�� ��Mn5��J�R'+��z̀w�U ��W ��� ��K���Z-���N��)	v+��Ycm[����<D�w���{�����ߟ�>Ӈ]U 4�9͋�^s`~~v�ͼXDvG�
A�yF;^��ݘ��j��۵`{�����@���A$qJ�� ���,��łK�h䘡kQm�)��B``���B��SI�MAh	�fb����7�� �r� �Ż���k��*�IUJ�R_���1�lX�.���2�����&n����>q`|���KfO�;�-X�v�����~�Քj��3�'g;a�Tu.{X�zf�CS�i���iL���N#-r&*��,������X�v���7�\��7'~� ϐ}�D���LJ*�Mp�Y�� ��@*�+�{���Y�䴊4�r�wq`�;� �����2{�ki�5���R�����]�p�Y�߱�~ʱ�� ��V�J�(x�>��8"��U?�}�Λ�{�	�2�ƛ[�D'�Wq\��d���N���͍JZ�Y%,�/;e��/w`�̦�"�W]:�5r�C�q�b��执�VMp�Y�� ��`��f��e�;!�Aj�|�X��ŀ�������Ĺŧ9!���?�k��7
��j�=��� �~�����<�`cyj�;��]/���� ��\��d�X���׀��i�쨎"�0�Y��f@;Ϫ�Ux� ~���"1D&Z�aD�����5��ֵ� N�i�%u��Z��f�pH YNiaZ��i����LWh�5�h�ۍu!A�-�vW@��3�%���=�q��s�8����N:;Υ�H���2ٮ�h�5٭�\�L�+�P�H�ncO��l�xI�#jZؓ�?Awƛr��u�+��t[u`z�}S!�g��gb�rJf��įjl�s�Y�p����mԫ]uQ;1Qlz�1�n�s'm��bu��o):���|}���)���f������||�k�G%�Q�+�h����1`�;��p�9����;�-Xڬ���RD��l*�;�w^ys��<������X� �6�`ƛ[�D'�U�׬�� ��@
j�_�U1*j4T�j�K�r}��V�m���u����=����޶FH��i������j��s�~���F3&����X��ܮ9UdeV9c�V�qXʣ�y�%S�$l[��8�8���p�-ݩ<Y�L����yڠ^+�z�ŀo{���N���'Y*���+�O��ϳz4D���W('�y5���f�ݖ��<�7D(�4� [!f�{���w��8��{� ����ߴ��Y�䴊4�r�{�j��e��?l7�����71V��
�l*�;�n���������ŀo{��~��+r��9��T�4Z��*��us�ĺ��B<tQ HЈ�:��w�c���wf�wf@-�2��P
��V���h�x�`�u�=m� ���s�@*���K�Z��UGѧ�UL�3�HD�T��������=�>���Ab�!6N,� o_�o7$��~ٹ'/ݚ�\h��T�V��׀k�ݘ�� �� >��h�{�&��j,ý�\�8�����3Z�=��x�\K{�jOX���ۅ(�t^y��햸��kx�#:���dK��J�׽��U��J��DĢ�T��n���P��@9vZ��*Md���5�x��� ��d��P]���ِޫ�H"�©[#r���׀u�-p�� �̀w<9�s4���AQa����bݛۻj��nՁ�V�X�ڀ��~�_c��{��ȥl�J�U� �wq`�̀w>�˲� �Xjz޽�t0'A�[Mni����!�Ӭf�,m�6�	*���#�c�	j�?nِ��@9vZ�[f@>W��-�:�m� �gu�ٯW�0���`�w }Ӫm$��*���k�9vZ�[f@=m� �}T �`u�bx��4��=p�� �̀w�����ـ~����G-,R'+��[f@;Ϫ�r��>�f@.N�{�O��ڀ �`kkW-�n�m�)I� ���4������W7!�٠��Uغ�H�p�61�U�D8�v��� g��l��H��Gk����*4TG$k<	Gm�L���\����/QE<8���y�
bs�V��@���p;q�zS;��R��1��q�y��kլ��gh�ɹ5�}��b-j�d�I%e�+\��X���K��˽�ZW%nX�d���G��sN2��l�ʺtrZ�V5�M�r\�6�r,*�n7i�;�=�x_V��>��,��� ����"��(�+�=M��s�q�ٕ���Ϝ^...D��O�Jӑ:�U� ���,�����.�\�`Ѭ�UR���/w��9͋���������w�0�&��z@;Ϫ�r��>�f@=n���эbN�a�p�]t6:�n�5�[a,��T �Դ-�Bّ�5�g�[XJ���n�z�t�s�@��ܠ�u�XD�7d����Ř�B�9Ç�0�������W������훁������� ��Mn5��ZX�NX�V�v�v|�Ϲȇ���Ձ��69X8U
�nU�����U�� ��� �l�y�\˘i13� ���=c�����t��XN��>��B�$���hYc�{WG8�u��m竞8��+s�Щ�C6w��]�,_�=X�ū�\��d�� ��x_tـk�n�#�e�4Bڠm� �>�˩\��d�kw�XjI��n�����.�p� �_p�GSp��W��lX@�<��8f�F��1`�})��D�\%�0� ��ȼ<Sa�G7�9���	D�<p�t5Ѥօ������A��1�HB0�dI+��1�%�� ��m��^ �X���0����y�h�[�� Ͼ�#	"i�GF
Gd<��Q��&�LI�Sr\epW���o����Ъ�B�B��vx_�Xl��,�z
>/§��v ��G�U>AH��!��x��D`��<T*[�G���V��V�R�PEr�f�����qC��M��yj��nՁ��U =�tX�-z�<5�k�}z̀u�d���.�p�u6ڸh&���<���!R�.�ݮ(�jbI�r��t	ב�<�0����mڰ=����9�}��nm�s(��AW�P���XN��:�����d�� �s.a�M���� �Ԯ��2�ِ����U��<�X7�V��׬�[fI'�g�]��1Y�b0nE��q5�św���wm�Ƣ%��$��`y�j��o;͎���l�n�,��[ۮz�u����Ke�K',�#F��9�N�v��h�6+!3ّ�*n���T+m_�7� ��0ͻY�$������jr�Q%W57���˩\�l�[f@;�W�K��6��4�vX2"�0�e�ͻV}��S9��Fi�`w���Y�奊D咬��� �gu����[f@/v�����f�5&�܀w>��ܮ��d�� {���ޞ�w�����o�� v�`˛�sk�[j��  ���V�E��'��+6gv6a�P��!w.5!��\pWPk����M&��%,p�0s�h�ݭG�TʭR�x+j�q�ܮr�=�Nf^p�8
���ۨ�(�.y{ZA��A��C���kY;@�y�b޲m�}q�׵Ӟz0G.ܑ��Ý]C�ɭĸ�pF���<ֻ{����UZt��Wa��qsk��و�Ӑ�1ڄ맸n���<Ÿe����]�ȥ�����,��nՁ�ݯ��IvC2s^ x7�Φ�%�ȝh�Y�}���6�X��Ł�m9���%g�3&�dj"YX��}�b�;��x{��o_��0���`=�57T#�q�+m+ޟ8�=�6�ݫ��'7w��;��R'
�-���ul�>�̀u�d��P�jo��Rjsv�����|s�$�9ԛ&I�˥�l�Мv:ɲ�l�#-��i��dE�+>���V�v�z|��$�����&���Ȉ�r9*�H��U�wwqe�|�@�`'a�)�*��ϳ�����OL��ŀo�׭���p���iX�ý��ٜ�\�&}�����X{�jE#R;�6�_tـ}m� �l�.����ŏ�x�a�k�}m� �l�.�������a�)hRY-,�V�%"!��m��R���)ѮJ���h�J�Zι,7�Jdx=z�c��[f@9wW �ԯ�����{ذޞ��vv:�m� ��\�R��ِ�̀q��"p��+��k�:�����Ňo�0�d!��� �"1�	�BF! *Xa D�@�A�$, �B$HH��$��ٙ����&@*�\ �`u�by��K�5�>�̀u�d�up?�����w�<�k9r��NY*�:۵`o�����nՀ��2G˹�]**8�{vb%F�c`n�cO[��ڷ�$m&�j2�,U%�S���]��9u+�}m� �l�sìԋQ��6�_tٟ�I&���Z�fZ�=����D<�P�Q�+Zv�`��b�;����8���<���y�������l�5,�
�`y�j��{�lG���_#�\8sMP� BR%����{��n�퇐��J�l� ��v`����̀^�2�Z�I�s�m�j��f!�����Ԗ����z���R\]�����ʥ�N�rYm���}l�� wW :�[���d��d����şɳ۾ŀy��`�����5��r9eq6��U�ou� ���W���̀_v�4謂�B�Ձ��I�n�`~�� }nՆ$�cy�X�S���'�U��� �̀U�\�ww�����׿������ +2��r��u�� _�]������Oa�$;V�t�M�Hu��m��9�n����K�9x�45��lZ
�O#�k����`�z�M�����I�ib��ӟE�|�WY%wD�D�ûf�о���Q	��m'e�n8�:p��8���@� k�\�j�����3��hEy�mm�3`��r �xw��^�Z�^�s��qq,�S+V��q�D��>;��+@���Z!�.�K�Y�&k�SX�,GHMT��QP��S�7����;V�{f�������8�C��B�Հ^�2Wup
�r��� Z����rJ�l� ����5�ճ��߻�b�=��X��Si�y\�j�l1$�d�M��̵`?yڰ��@��kz�ǆ��\�ِ�f@/>�W�W M�Oc��cs{iW6vڻ.����'k��_w�ܜ�e�����+5:�'^Fa���ͷ����� ���^�\�ِ��F�����2j�.�nI����uE�!��U�+�}�f@/u� ������h��@*����̀^�2zw^ hwu֢%�KS��0?���{3�1��`?O�X:ӛ�F�aG$D��B�Հo{��%���}���7��,���W��YU�XG@�V㗜Y�6��nQu�p��b��;7�.�Z�@vu8�N[*�5��0�l�_[2{���;��y�������U��/�� ��d���\tX�kz�ǆ��\�ِ����O�`�*�F�R1!�B�,@�x��*��/<�nI���� ��Rj4��hXn�� ��d���z�p�f@/�U{�1n3R��
���U��/�� �����uͥu�[�ȥvA��q��r�Q��YL�;@���;k�"�1+d�5ݦ�1o�O\�\�}l�� �ݘ���Z���-N�J��7�ڼJ ��Ձ�^E��9�dn����z���@/u� ���^�\�ِ�[pŬ�n&��{�U�$��t�,�bɰ[�a<IRK�2$��,��vHBnD�#$��x��!,�*B �h)ϳ϶nI<�|gưƨ;�����l�=���/���`��xm�iͭ�
9A�e^�Zt�+��n�K1:)o[�l�Ԥ�.��$���6��l�c�Zy�}l�� wW ��+�{ԩ5i�B�u�V����.s�\�2ɰ2=�&�}n�yqq6{�_��H'T+`�X�_� ��+�_[2zِ
�90֖1o���]r��� ���q$��� x;�:�D��ju�R��[�`N..,y�]!�P��{7$�
 ���U��
 ���U��
���*��
 ���U�dQ C��P��DV�X",Db*  ��P`*@b��Q`*@ *D�"�X��  ���"*� *(�`*�"�(�X
�U",X�,T� ��F(��"�@ *U"���"��"�(� 
�T",(�X",b��P�"�",(� ��H",F(��"�"���", (�P�"�  ��b��`
�X�,",��*E",E(��"�@"
�D",",b
�@`��D�*R� �*X",B �A"��b�QDO���*�� U�U�(�Q@^ �
���*��
 ���(����
���*��U�U��
�2����������?�����������}ڂ`kf�*�@ ��        � a�R]� ��B�iB�Z��ۡ�5��euӢ� � "t���iqe�%6eŔWiGݤU�.,��lzw@o  {��浒Y��(���ጥp]ִ��$�ٓ�ݛmol�7� $9��@(��(�P
s�e' ]қ�9v҇	�J�  =z���T�ceWy��Q�sP��� �@ d$�IC 	� M4�L ��UJ#J�0 �`  F0�2d�L&F@��M#4i���)R�#&db ѓ114aB�4a�M	��$Ѧ	�M=4�)B�Q�`  ���&  ػ���u�	�� !3s��QU@�~�2��� Q�D
��|>��*�1~����������$�+������͟�Nؾ�=�c��m+h�ߕd' ��m���ֶ��¨[M?|�U@�ʕ�o�I4Q5�c=1r�Et҄6��!U�XJ���2����;�[���D�M�DU@��Ɨ��cN;浃��[Z���?S��!�>٥HL_S��&���D�ޛ]w.ִ��)�>3�{�|4zɕ����Mzx3DX���b��@��r��f�0'(i>x=�`x�[�<J-wF� �f/+j1�F�&)�/�]�T�I���ŕ
7[ޔ�B2G|��A���".â3��`l�W���`"(ۍ�"����mE��(�Sƣi�i3*�`&!@��D�pu�������$ƃCh
�� �d��`7I�`"�n����D�A���#c1�An���t��!��u����Q��[!��i�r�;f,cE�tw�t��[#dt��H,�N˧s�6C����z��-��:Te޻�V�QXYXc䙣+<7!`Zn�1�]�ZZ�wni�����
#��`��\��dŔs�s�(��� Ƥ`���;&�A��k�P߆�khS<6 B�Tڹ��[f�w^��!>�s�h\��1��~���:<�s��i��3M8� ����#��@vwf���iVl�Iiq�Ŧ6�!������ǀgnB�����ޜ� �����mp�����A��a������N�"���Yl���v��k6��L1XZ*6rc��u�r;<H���Ȋ����c��>%�ղ����ʍ�˼�[�l&�oi]3����[yē��Tl$�xa�wפ��	ӠݮD�ND��r:A��#Ll�:����;<b23Q��d��-�&kb8�"&�k�ŵ����$O��[☀I�6�6�Q�y��1���tϜ�<��Vd�-���`��U��W�@�$t�Ɩ].wF��(�#Ѽk���H5�[�8cZ-1W0�f���ʴh���/$��d/"�01юal3��0͐Bo�C��	��~/UU		i��������%��n�ok�J�
�x�z)N��&SȄ�5��4>hk�Kh�'�Ɗ�1�Z�HZB�@5uP�\��a��nr�|�C�{Q���#sA^\���48u�"���I
�����ǋZ�-�X�3�,�M�%Ќ���}�9����>g+�WlkF�dG�Yc�h��Bw<#Q���Q�
��$Q�Y�A�-����#})��#{�V�x�{Ԩ|�M��'8OX'��k|�l�ʉ#vO61�ㆊ�qz�	��pyջ���ӹF�0�i8h*z1��e-݈��d��#�N%�w}��LѲ�8w����0�4�v��&)#y��q:�9з��ӳ�Ն�j���Ѡ��#�6�Dhb�p�č���:h ��3�㰞��ZK����0b-V��׮&`j���1dlvq:�`��쉱mNݤp��F�%"R�T��tI&�y�|���D�'׆|�Ǒ�3v)mZ�pB9�j�G6m<x �-gT�A���I�7�7!v�놃�������f{��EZ��O�yc7(���#��$��wf�͐��7M���ʵ������j�T�V
e��O��W_���}6]92�̡�RP��c\UU6�W/]j��1�'I����a������)�U/�RŚ^\d����;�w�y�$`Ue�j�SCWlR�oM�D8��⬣P �WZ��.0��=��f��E-S��(4�Y]���xXe^j��p/9�W�:;[Q�!��k����L����;m8ܔ�����/O�fvv@'7I6�$�ԳbѪ�\�&y��ϸ٬c�`�c/.]:W$<�kH���-�i7&�����"@�m�X[X���FtUUV�t�n
����u�;"���ۣ��Ph�ƫE,#��.����tn�H���)�^�j�eJrc��*UUvӖ7M��q�|�u(����^jwl
��@#d#m�-��^4�a-��lj1q���ȤUi7��
�X�r٩v��ݱ��@N�+5ʫ�Q�9��u�Knin�v�yY_%����
^X��VtK�!+;����U*��pյ��%�S��j�w��i�X6鄠jt]W['��[|�U)6���uR�sUK��Ok	T����=��Ί��I� -����K�R�p�B
Y]�*^USS�5Ur�Sf��j�6��V�PdT�W�	�s�JA�I,����� �K���r�UK�t���&wh�M��r= ڦ�U�q�z�R[Q[L�jی��9+'U�R͋�ew;]uA��QӜ����v �;S]J�����|�ʅ檩
K�r���Ȳ��[s ����A��8������E�5��uU*�[(�r��W�5U<ܬ��P�s���rUZ�D��୚g;X�X�u�W*�T���:l͵	��������ψwσ�-Ǫ�e�$<�N[kj��%J��J�� <9���l���<�m�]e9mUU*�*mWt�[E�@fʲp�IN�=��s�J��2��UQqe���V�<�:�vR�;Pq/��%Z�Km���wc`�[pK�Gm���&yd�P��*����D�)[�
z^�!+���Ͱ.S#[H	ҹ�/.6��
:�p���Ƒ�o.\� n�\�m�u��AN&Gȼl����!�J��WP����Ī�5MT�.^����N�JN��� 6`R���B�nh�u��V����V�._ ����E �ѡZ�V���km�VԬ��jV�d.�he��ـ���j��UUUX�U]UuSʜ��^��V�UWK��f���MS�v��U��n��  J�U@UWU[RNMMT�����v�U���i2g�`v�9Z��(��U[l��������W8�%��YyyY�Q�����&�j�k�.GN[���'f@���N�֍J�ղ�[5M/2�\<� ���i�ڙl:r�n8)����JEi�Z�X���l��\M���wW* <���u�����A��Ǥ�����}���� s�3ޭ�aXD����B²qZQL��M�h�A@EI�C�q҈���"�l8��AR������Jx����DI�>
����SJȭ*x���h�S#�Ya��Dq�%�T�x�tLI×Gb��؋�E<M�j�Y����PRBK�� �����lTe�TBj�n��IGj ���A�FE=�[I���_8���P�J�:�P!�!��P�s+Ԓ��g��4Z4H�8T�k�mf�H��m�N^x���e�ٖ�8��ՋNQ�c�n��������M�6���ӽ]��6z葧�N�f�\;t�_C��;�!���g<q�Óy�v�������wa���n3r�=^L�v��sk�G!�J�6���:�w �	;ay��W=�۔�ʡu�T��9��/b��Mc��5ی����ǧgjN��)���d�]Lje����n�Ǎ4G]�83"�ex��B޸,���8���I�nNF���ժ�4u'	l/%:�ZMk&�R���	��[J�Vh�&����pN#�k��Y��-s/���]���\ok��������Z�����oe��Ժ�+� ��e.n%��&5$�F�R��?����'$�N���~��w�i<.�=��e��|���%!()�5T�Ф�J�*�E}����Rl��DD76����� Npt�wk�+�rKt��)p��
ձ�̡���W�s��|��)˦���IM�K������w�i��sZ�f��$��D�J�[am����e=-�;௓�[�nfNx�R�nl A��M�wM�C�K��%	biI�UR����2���{���[����M�]7v��K���(���o�os ���bK�a�9�E�QZ�+E�}���\:�Ŵd��
���E�9�-�{��ЙwW���弶����#{�|�r��GEZ��t\1;|��_�>7��I�������.�>��2�c��n���sZ�m��*���[v�pr��Y55 �n�I�� 
 	���(���n��|���;����  Fn�qyF>OT�:�A�[��i�]�^�)�<�������^���[�v[�R}�pշd-�ĤQ5TffQPd�J�P��n��|���;�������ۢ��FL��)��}��U	d�K,j܍�]$���k�מW�~�{��O�;[vQ���n��+]2�n�Z��i��e*q�p�ȘƇTV�.���O�|qզ3����F�qD\�Ӯ*�I��m�6��&�/�v�������$�h�������GU����Z��=r��n��w)��}�� ��w�NZ�/����zH;!
�m�W���\��c���@��@ �  8󕮙�[�ws�8Rv�������w�+�Tȑ#��-�%B��T��|מM���޶�����H�� ������\`����w��'�m�,�Q�s M2D��!���f��
�X��HNY&6 |AgM&\7ú21q���j��V� �P�d�C#����
�.^)-c�6����wk6���R�:���$��DWd��/5�O6�U�ۻ�7n��n��R�c��Q0"1�`@}SY$-�w{<ܩ)*�&�����WE#%������4~_ll�vQ�3��c�V�K	�ww=��'���`D�@1�o�����<P�G7���>��~mQ��ٸ��k����7p�k���ˡ�i�������v��Y,��ߙ�;��E�������II	-5o�h�����}��[�w�E�K���I�p����ßkL����X@Nج��`�����~���^j����&�Y�=�����+ov�J�6ݝ�.N;�gN&��7'�������v�>s��{��:4������$��ë1 AnJ=�|���畣�b[�wc�/		�j���"��A
U"���2,�j,��tl3j�!oIrfQ�c����1d22@� Y�oY����(�j,��fQ�d��IԪI,�X������"w�Pڌ0ȳ� �V#�7b��hI�	Fa�<" ���64�Z��~���2@`݈R�%�E:*�u��\%V=�.�����Qd2�&��5��n����-=��]<�����o}����M�j
�-�\��XL�o6g�0�}{����C1v�z�I�E胺�)'��X���!�'�Cj0��<��I��QUd���U*���h��1D3hm.b�g�"
軧�q���o��8y;�z��{=��IZ&7Ta�E�����!��C��o�ݛ� W��y�C��������1�&���cO�cQ�0�O�O⡵B2,ǦѿR��b�f.�ї=g�-<�^lȼ�=V"Gehcv�)T��Xf+3B��LL6�2,�uc��1d3ho\�)dQ��� ��93d��,i��Ő�LJI��BX��Y+O9Ǜ3�ўM3�Jn�!��CF_T�a�FQf6O<J�1X���t���hz1�a�]�)�r�ۨ�t�^l��[�rŌ�I�����p��}n�9ކ�L�0Faci�]�a��\Č�f��	�1�Hİēse�q�� �3n�!� �:h�sZ���0�1,3B#,
��	�\0,Čs�8���b�$�F!���)*�}3(�.������"#f�ژ9mE��3JC,`��vz����m������T�ϧq�;����lګ񭩸/�2pq�ځa�^�[F�t�n���� '���u紼���`h-�I��y*�ܺ�p�]���܆X�U2�4h�܋ZE�&y���\CF�#n�-X�ڡ��X���+�^��wj���s�Tw[q�<��:"�V���J|(�Y�v�k!�MD��Z���5��:{l�"�"�ۑ;B���8����2q2��ٷ\�v���y�2q��$*��$�5�dY�,3���b%�_,J%���ı{�zW<�e����js�N��^yP��i8W��=�[���&r�7؄�qָxuqPn"����R����<K��묊6�n�rT)YZ��'����p]7���qv6gEFQf�~���ő�Q�m*7Vp΋�f�}v�}\�t�.�5��6�%�Ik��t����0�
��<ѝ��qM�� ��1��� ��I\&7Ta�"�}��$+�b�f.�޹fJ0ȣ����}�O�.'�.�壶�O;���;��}�O���<�O�V3Ҧ� QE�	1v���`�ȣ�d�\2l3�2����*dH2$d�<r�Yp�uL�ؗ=kfy��B��!��C�r�"����@ֻ�~�����0�q�@z���%��",��߶�1� 2,�m	*]I+B�B7b0�X���f��UgREm l�Iɰ�N(f,��%1#�����0�z��
ᘲ��<�33|ߴlV��"��5B�潎�M��5��V���v�hv􇡻���E��k�߭7��n��=�6PV�R8_�i�F�oT�3�S=�ԲfȪ���b�C1d"yy�a�E��63�M�1D3hh��L2(�j,���"�*�E	T��~����mt˶�zGc_~��M>���>F�[�!\i�,}�6����%�(�hh;2ݿ��K�|��3�l[��G$���n֤�G,�q�8�fs����]�}�i�,�1���$�"LD��C1s��&��F�L^��0,���+D����l����@�����a�V�.f�HYb��hw�Y��3���Xc�C7 T��H��/i�!��<-��>�N�<۳�Ϲ�gLиf�ו�SO�%��,�卻d�1U-�:(g{ՙļ�~�M.�6� Y�}�;&cu1�<F���HV>��#H� �!�t�@ia�,����v���ss���Aܕ�ěf�٭u$���#��W=�.��0�l>ܾ�4�j�We��Z�^Qn��edq8:���{��=j./��薄�������D@�i�f�
cW�li��hxgب��"�n�b1�׃�]2m�	hK�����NQX�m�-S&��6�cz�8V�"�@�(Đ�e!�r̤"���;�ag�"Ƙ�A�� "I���a�f{�꓉��!��V(�Ub����C1v���TH�0�@���&Ýw#�x�!L�N��;�(	��͸��������ݞ��zm��s���[���A�e�kN$�0	�I2��Oc0><3�[��=$�m�zz�g�`�ON�uH/��i�$���?G]y���ui�v"�}Չ°�C1v��j��(��5TR�Z\�����*g9�bK�������,q��΃$�}��u ic�lb���4� ��!)!���%.���S<�	o1_�3�+r9an;L���X�c�N!�#�S�0�@dY��8��d>Lf!޹�H��Q��ш
�^^64���d����4Rm�I8
��WBE�U������v���7j�{��6��燬�Gu{L��O^��Ke�H˓�1%�3��Ӫ6�u�	Q,r�J�ǜ�[�g�im�4�����UK�߽��y�#p{����a����YFc�F;z�*F(ڐn�2�����������dw�\�@fs�a�aȡ w}"����D��p�p>�d#x����/���l[���9(�mܲ��m���%�C7�ք�ޟ���6.	Qy�sty�hɘ��3;�<�X���,��NJD!�E�dYd�礍�d���VE,�7]4�f��v ,�'�.2,��Q`#k���l�gq�������n|�*b��G���k�*�1�!��#�$���IR��h��Um�G���ōh�z״�@��?����H��Q�"�6��6< j�F�,�O�90�\��,��疻MWr�݈ln���J�qJm���W/�ւ��s�b�ͻjV틴޺��9`�9���g�%uT+[tM�X�U�k�ZODY�(�c�@#�M�1�ΐ,��L�2> �@�d#}�_p4�%�Ŷ�f���p���P%��K�R�:ެlK��s���З�~����G��󆣐r2��׌�9?���c����@� d|>yE"�Q/5��d�-�v��IG��k�l]���&�3g�1�?~o>�\<����3��cS4b� D�L2;�=)c�M��^��,�]е묎H8��d(���e`;rfš-�,kFv�z��K�Z�Vb�队˟r�4�(gED��~���3Q���9�rr�:ژֳG.%�Ĺ�c����l}��!e��i���V��.E��n6%�Ջ�8.AϹ����%������:F �QՃ��U� tDbb�C���$K$0A󄩴S�����K�����Ls1�	 ��`���N�s�&��t���XNf&&�E5���IAc�c��΅�S���0�a�T�5K$��0��$ԓ��Пټ�;�F�8"и�J>h��$&&�nΘ���nۆ��赝���'*zF�
�-��]v� v��n:�ä���m��]X'd4���	��9ڸ��q��45�^��U��<-Ry8��y�.]�`d��sa�
$���<GAMƶ�<�5ݝD��I��s�
�E����1j���d��ӘBm��"�m�q�.n�N6Iz���R����8��gY3����:�)[.*]2�Z�m�譍�lL�=ewF�Sî��Q�\�z�1�����%�L�&�ka�����kJI4�t��� r.�Ads� ~� ?>��oY͛�f������e���47F�m/��h��P^�kn��Yk;��³�+�n*���s�%�l�*���^ވ>F��Ep�w����g���'{읪Sb�ic�R�1c� 1�t��n�3b�l�e�ץ=��l,"#���#��I�J�M���:e�v���S�=�舟U<;:�'�k��u�3Gs:f��ߺV�3fR:m{�l3� 5b�%�%)����"�26��ٚ3|Y�h�|��uk:<�'q�����Ocq�$
�(� %����'��^�5�\?)�'��!lP~�L�3b�y��$�hqT�u��V�Ҷ���8f���IB�o��2|�Ogw�D>��������;����������|�~�W�u������e��e�dc��Z۬����b����2(�1F6lt�l3���Bc�a��E�0�1�~+�5���������a��9�a�9�/4�y�i]� �V���mi�ϩΊ���۰v]�A�kg��]tO�j[�Z�Q;�J���,Ėz�?$��ǽ�9*��*˂r�*�WLؼ�f ^!�����O���>�_�0@�=�2Q�@/P�F:lzX����b�K�iE���:�u(ܡH�EM0ȲhY���_T�d`�
��3P�G���H 6����aӋ�cLa�v���d�2=���3}wԫ���G�<��;qU��-��F��ڢ��c�����G����:x����?w�$~�~#�Xm��?%�]��uLط��nJ)(Ipb���+dis�S8-	y5��M�~>�CH�hx��rjc`����Ӈ�w�yQ� v�p""��ڢ���b�#�dmY-`ծ�Im jʦ�ٜ3ZBA�0�� D���EW�}57bi1d|2������Wr�f=6��M.��Ş�˞�޵�x5'�l�����"�"����9,�՞tN���Buո[���ƹ���g�n�`�wiH�S�ӇZ���55Ęm1��~\3�#���;��#����#�f�1����͏@�P�i��$��Řm1~�bJ��j2�)m#�Y��Z�o:d�t�X-��rY�X�%Tѐ�}����͢�1�4�ڎ�,SC� �\cw%�=����p���}>�$ly#��S��Y��ēԳx��ƴg�h�f�ܤ��a�b�x4��b�c��('3M$(��2F���5�Z����`��`�&$ ��X���ŧ``8~;����B� bL,�YXX��$�c��HL������$�$,����|��I��&��Br�q ��h။i� ��0,� �fJf��f �I���%� �0
�dd��Y����d�(��(h��mG��ju��/��?'V�#� 8GQs+Ҍn��(�b�{>�Qv*�T��R�c���t͙���C<�E�F���f:�x1p�f/��c�����>��'��mM#1$�>Sa��@�C<�S*fa�8ҩ��67(�pZ�ю��V����=%ɟ)�,�� t� z~{D+|tƑ�г���ਗ8֌�ť�9Ϩ�W[����u-^�7e�}�f�s��j�5�I��Sb�.�Z#%�m8�A�K��\KYԖ�m��7`�-�ci��K�wA��bb��S����1�a@z���M�1�i�	$��0Ȳhx��S�/k���\3B�?`��ae���q�@t�Ĺƴg=Y�kb^_=��(`�	�t��U�1�|" ��f=T��lq1b���sAk��_%�,���-��B}��X@NPluج�ip͋��{j���D�o��]��p���~�p�w?lЈ�t͋�j�3�#ε�:-�{��(��и%�5�H^�c���N��(�l��bIf�*չ��<kF{k�qk8fbş@��޽��cu1�,�M��)��=���8qO�y�Z�R�E�
��&�Ɠ����;[�_��p]ř���ε��h�����8䨶&�����p�ָ|��}NB}!��?�v}��#��{����|�9�/�ӻ��T�������}<8�<�O#��}�<g��\!kK�c�$�{O�%�$p&+l�^;jKX�[���Z-ў8,�s5���+��S�c�X
z�31jW�`gz֌�3ɳ���p�{>O9���5�F>O#����܃12~ߍv���>��g�����ŷ�3f}�>t�Hڮ����),���ќ>���g˖�G�{V���TN��|������'��׳�}�-�$`��[�3a�����M�sfp�i��9vD��N+#D�zތ|�O�~�l�w�����~N��о��>��q�
b_E�S3�5�T���bLo���b�3h_�|2�1�15Y�7��À"�3��+4��҉"�J��9Cy�7��f�������4�#� �S?)��0� ]�$���� 6�.��m�FƐ������[���'!KP�f�@m0Ȳv�6�!�.нG�UC"L|wP��^�l}���G�Vy���0�����D��1��{��Mu����x`�D�0���9��d쬈�\-�W�hNl�y�Fb���.��������F��:�7�����9ڸ�M��o@�k=������[��m<���{lv��M�Z��bȁ9U.89[��P�t���ݝ;���I�We��Ν�ϳ��ړm61ʀ=�=8��8�(�X�,��0�a��b9k;���s�RŬ��8���ݮ��5v���=!g�;��;3�6��H0���;m��R�{m]ѰIu�n�v9�q���q5��n9չЦ΍ֶm�[!p�KL��d��7j����*܎I-�[.��x�x�f.g����(�x���Z��~�6�RI"�R+T�KF�lk��۩�q6�rm�sv�1���j�^��E�f��b���������{��~{���e˧��uQ����1�2>#1
'/�"��g��>�E@�_1�}%���@�B�2,���5ƍ.E�-i��l��'h�$-�9J���A.s��Ŋ-����p�%���F�6���0��>��{�г� l����h|)�^9�(JOd�J�`�%'��j��`�%'~s�k3F}��ֲ+5�Z�5Vov�'a(Op�(JM���J��(JNɐ�'��n����(JO}��%	��(JOd�J�`���)?��拉�J�`�%'$�)�H��P�����q5	Bs�Ǜ���I�L��.X%	I��&�(:>k�)?w���q;	B_,����MBP��	BRvL��?o��#q�*�)X4R�Pib�����J��P��ɐ�%��)>o�k>�8���=�_��%'�d%	|�J��15	Bo/��Z��%'�d%	v�)��>bj��0J�[������%	|�J�~bj��0JC��x�7&I��'��ݮ�W�)=�P�'s�)=�!!b65� ����qv Z�RYk���3Z���'��P���!(K��);�MBP�������(JOd�J݂P�����J��P��y���q;	B^�%	I瘚��=����	B}����pJ��q5	Bw0J��2���	BR}��?k8���>f	BRy&BP��	BRw����9�v��r����[ֽ�r��n.�hxҕ�v������6_`�����!s��Z�f�n͞5�۟U��Ξ�R4��=���n�\�$�ơ!��"��Ո ��"�P�����J��P����϶�'a(K��)7�&�(Os�);&I�RL�������\����P�'s�)>I��%��)?~�.'a(Os�)9&BP��	BRw����;�����P��ɐ���s�	BR|���J��(JMn������dq��+L���kň#�	BRy�&�(Os�);&BP��s=�\����MG���!�>�!�5	�`�%&��J������=�����v���%	I�	B_,���q5	Bo.�u�Y�(JOd�J�P�����J��P������'a(K��)w�&�(Os X��LX�b��`��T�P���R�t�CK,A��x��N�	BR{&BP�l���y��踝��=����	B^�%	I��j��'�M~=޸%	I�L��-�%2�중�j��p��|���J��P��������%C�J��q5	B|����L��?nן���%'��j��0J��2��5� �����)>c��\�-���e��޳zΧ��'��(JO$�J�`|����MBP�����k8%	I�L�`N�>��=��%&�}�����J��(JM���J��(JNɐ�'���W�\����MBP�����L����U<C�lL�P��O|�.'a(Os�)9&BP��Q�1oo X�ƽ���s�!�27�9��{�D�)>I��&��(JO�15	I�w�������Ǟa�#�S�@6�dY��W�Xf0�c���KOң��hY���9(�T(����� �V�4��n7]����@x��89/n�̻������]%����rn�^8阮�������z���Sk�Smp��{��K�|��C#��w��cLQ@�B��ʘdI�?�b��_c��3G�~.�%(N�E$�D��ѥ�5�8-	vo'�M�S"����Z� ,|����$����R}�6>�44�ؙ�����5���ؖ���hs��AYD�n�q�Kb4�e3�kMk��[�8d3�a����>���sӱ��j�R>>�s�jkaA4bXtc*���q��>�{�c�ӭ!����T`a��FQ`F$`�bNV&UI�e�a%�e�82�Tb��dŃa!c�Mv|�Ѡ�E�\�zA��5�C8y�iv�:(3E�`L�4�	C�f��3�#��j1�Fc�ac�AΜ$�}$�UM��T�&E�j P@�QPt]2�P�S��||UA�Ks����F5��8c��d��a��C�U���"n�2Qȉdh�۝2Ln�f��7�E44��SGҌ6��f,ǆz܃a�����,�+��u9�~,޵�=��:�$�� J� �
��*
��A��=%a�F^����ǧv~Rl3a��BM���SĘm�~|Ӿ_}�n��u�<�F�'x(&��o���xy��ƴr�qe �d��a˸�[[;���)��\mӬ4�I�I�׮k�tNE�3K3Ie����9Tu��L���f�֌�3ſ5��b�3k����cLI��,����U�1��1dt���0���6c�3�_o���#u��Ym�� �]3fvy�5\?k�����\)�Xr��Ü�ߍ�16�g�KG���u~�r�?��s��9��pNѻ�%�Ie��}9�����|>����� X&4@
 X���ܟ�} nn�L��K�n� [�鑸���"M��T�DX�{5� �8���w~�r���k�*smبz���y��v9�$�(R�&�#�JA�D�&��ͻ�̓�Nۻ�6:z]�v�ܞC����
�lۻ#��6�|um��Ļ���SE7nSU�{C�L�������s��t2L�lγmΌ�LM�K����5#ӶKi�*�!&jP�j�'8�����l�v�9�)��|�b��w��'�?ٻ��v���$�!b���H���\�<����D@�!@Q���	�})�w~����k�U:�죩%3�$�T�RQT�Ԕ�c�X��&�����Z>��#�!: FmI�����@ɓ�|�{�s}߯�}MYm��:���T�R��w�y!?�=���T�� �;��~�K�1�  ϑo��;���=I��9��\nIJ��s����7�-�n�7�����W�t����g�MZ�~y�g,DR�+��W�N���+��hU>j���^0��>�N�j��z핵��-����k�3�:���Mb)L�sQ��N5�$ޮ��ac���Q�]A�nռd��ny�&��ˮ��칍��|>m��<���g�5��ݏ�
���+u'�tq��grO�MX�b��s�Fŵ��g�iq�]�3r��<y�T�!������=r(�n���6u��p.p cۄ�K 7j杻n���q$v҈�zb��;D[#�ۄێ.�ݪ�Hsd���[��6�,����;u��A��Z�p�Gl��uv��퉤N9Q�yֈ���۞�v��U�ՙ���}�
J,�2�������A��}��B�Φy�P�h�R�`W��}�Q�ծ�3qs�GC�˃��p�*�Ud�ꔑ��)ˋŋ3�Y�hǨ��ډ���d,��jk���o�)��|�g ��v��amݩ7ǩ?�33�{���}�k�n*�pC�q�R����3��^�;���y�9�[On���]�v�s�����T�L�Bf�*�2��5)UJ-�]�0����U߷��ր�JA�.!
4D���I$�Q���1�H@" ���ܒ9�L���B�]"[�����nE�)#j��$r�^^;��{˻n��p�o1�+Yҋx�@���qS��ziW�޾w:e�<��]��B;#���d����W۝����ϥ|wr��Y��%��73��&�m7w>�3)ݷdH�6ĪT��ڥ:��[�#�b�V�WzSOA�pF��a�H%�9l�M��n�`Ȼ�{k7VL�nñz�V�j-�;�o� ���;��m�̞�.�H��ſ !����	*d-
��VB��c�Ns\ֽ��ܥ���
ws���w~7qt�	[�����h��r��<�	�FW5K,�A��;���Ƌ�n�6�ro2lP�y�U.�:���e�ѧ聏s.:�)���2+jr:�r7(��n��?7}Ro��/�rZ%�wk��%'m�� ���ҝ��5����M��d��
�[*
��ǘ�B�]2[�wٗ�F��w�\Vݭ��2�c� hg�Δ�&���*�W_Kk��mgX\�jE�Ƽ��[�KЀm9����"���z�m�:�@66��of�OWNF6�[	j?Db4SNM {���x�	v���M~4u^�my7��B�]2[�w�K��$�T�"&X�"VӖYK�s�ג��N���K�c���xL��w�NKD� ���^�l�ֵ�ԍ�$�܌�:���IK)Nj[���ܛ�w�f.�-�2"#{� �:O|ә1��#�iXH�W ��6��R�� .-ȢdbB���%���̕-�u��e��]m��k��um�G�Hr$ah�T�U)�-�?��΢wmݯx�$�n�gVq��[���PDA �ד�����{��D�-n�s,4ʩݿ� �̵���@������;�y��gw1߽8�"ݻ�"�>���4��sz�� t�{pg��n.����받� �ѭ7l���SM!pgUmsp�%�{k�����n�1X����k|�7�O9�N�s����ӻ���f/H���e��U���C��9dq�rIj��vZr��s�{�3���`���ߥ�$[�v��2K���N�R�!o&%"���P2f&h��"������_�d-�wuu����<�,U,PL`�᫽����6ݭγ2߃{�����(�*d!5T�55@��3T�n����2K�f�e�DU��s�i�-�?D &�@ �!��ru;��ZRT�r�)4%L��QQSJ��m��R�Eͷks�̷��[�v�d���'~���>�L��nv㛋������u�x7]m=�n�v)���􉝼+�Y�s�W=��
�ұs#ME��!$ecVG��Kh���i�K���2��Vy�-ۻ��<z77s;֭�wM�ٻ�di��M9Tv+jr����۾��(�؈ A���2K�wjus���#cg���u�xI���3BU
�T�JB�T�In��M��i�w{֭�w[" H7qUu����N1E7n隣��*������&6��_�σ�.��=TX���e��W�䟆�� tP`H�fx�i�f�g;�2<2�Х*U"���*R�.�^���o�ܡ�OE�{w�R�ItߠDDɮ^ڃ,��q����I��DA�$��DD{f���'ֈ��`I�OD$z':R�-��j�nSr���((%A܀:(�P>[%��N�x�<���?��RP<�$E��4G�^V��p���̗���i~� ���ǜ�Ō�4{���B0t�����$�fm'��q�#]���,�P/������+�yH���� \���~��UTj*��d�GqS-��k<�!��߅p}!ÞR���u����9�M&��p�"*�iN�5j�Q9��#�����ó�aV����IS&�KDdF�WՀ�=��~�T��[�c�˻���ө���N�M(���~P�GJT�ɪ��P����� �D��0
���� �A(� ���y���3�P�4;k��Z�E��b�~���(��Sx�sbl��1�[a��	������?�	���H#�p�#ăQi����{�B�EUP!6�$������k��!�N����H��o�N]���0�b�;��������������燄i�OY��#�����f�i�$ET{ Ą����y�&%q>��{��m>�]� �	x I؈���Q��(�\U���3��"�Ɍ!��b�U@�d�7D%�PP�������@h�y�?�ӣ��+�o�:w�M��氬�/x�?C���L�LFJ|���ΓZ�(���=���=Fo0�G]�;����q�5�3���N����Q=����������d��q��Ǖ�����5�4N��ɺ <C�]Ǧ�<�L}�Xٯ�P'_���ƃ�&�� ���Jq9i���DU@���8s��ӳ�s�v�e�����)�JC�x���li�\`c�qݽ*a�@�����1֘�n��N�T��R�~Y��4�*�W�P�:����b1�T�n��C��D^K����G2	���X_�p��D�>k	����   C��P�
��x�~�=�O�
r�dT�u��0��-B\�)�����0�Q�������B`��x�%��Y�3?���)���@